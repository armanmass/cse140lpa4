// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Jun 3 2019 04:04:58

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__23195;
    wire N__23194;
    wire N__23193;
    wire N__23186;
    wire N__23185;
    wire N__23184;
    wire N__23177;
    wire N__23176;
    wire N__23175;
    wire N__23168;
    wire N__23167;
    wire N__23166;
    wire N__23159;
    wire N__23158;
    wire N__23157;
    wire N__23150;
    wire N__23149;
    wire N__23148;
    wire N__23141;
    wire N__23140;
    wire N__23139;
    wire N__23132;
    wire N__23131;
    wire N__23130;
    wire N__23123;
    wire N__23122;
    wire N__23121;
    wire N__23114;
    wire N__23113;
    wire N__23112;
    wire N__23095;
    wire N__23094;
    wire N__23093;
    wire N__23092;
    wire N__23091;
    wire N__23090;
    wire N__23089;
    wire N__23088;
    wire N__23087;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23079;
    wire N__23078;
    wire N__23077;
    wire N__23076;
    wire N__23075;
    wire N__23074;
    wire N__23073;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23065;
    wire N__23064;
    wire N__23063;
    wire N__23062;
    wire N__23057;
    wire N__23054;
    wire N__23053;
    wire N__23052;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23031;
    wire N__23026;
    wire N__23023;
    wire N__23022;
    wire N__23021;
    wire N__23020;
    wire N__23019;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23011;
    wire N__23008;
    wire N__23003;
    wire N__23002;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22994;
    wire N__22993;
    wire N__22988;
    wire N__22985;
    wire N__22976;
    wire N__22971;
    wire N__22968;
    wire N__22961;
    wire N__22958;
    wire N__22957;
    wire N__22956;
    wire N__22955;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22920;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22891;
    wire N__22888;
    wire N__22881;
    wire N__22874;
    wire N__22871;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22849;
    wire N__22846;
    wire N__22835;
    wire N__22828;
    wire N__22817;
    wire N__22814;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22781;
    wire N__22780;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22768;
    wire N__22767;
    wire N__22766;
    wire N__22765;
    wire N__22764;
    wire N__22763;
    wire N__22762;
    wire N__22761;
    wire N__22758;
    wire N__22753;
    wire N__22748;
    wire N__22745;
    wire N__22744;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22724;
    wire N__22719;
    wire N__22716;
    wire N__22711;
    wire N__22708;
    wire N__22699;
    wire N__22698;
    wire N__22697;
    wire N__22696;
    wire N__22695;
    wire N__22694;
    wire N__22693;
    wire N__22692;
    wire N__22691;
    wire N__22690;
    wire N__22689;
    wire N__22688;
    wire N__22687;
    wire N__22686;
    wire N__22685;
    wire N__22684;
    wire N__22683;
    wire N__22682;
    wire N__22681;
    wire N__22680;
    wire N__22679;
    wire N__22678;
    wire N__22677;
    wire N__22676;
    wire N__22675;
    wire N__22674;
    wire N__22673;
    wire N__22672;
    wire N__22671;
    wire N__22670;
    wire N__22669;
    wire N__22668;
    wire N__22667;
    wire N__22666;
    wire N__22665;
    wire N__22664;
    wire N__22663;
    wire N__22662;
    wire N__22661;
    wire N__22660;
    wire N__22659;
    wire N__22658;
    wire N__22657;
    wire N__22656;
    wire N__22655;
    wire N__22654;
    wire N__22653;
    wire N__22652;
    wire N__22651;
    wire N__22650;
    wire N__22649;
    wire N__22648;
    wire N__22647;
    wire N__22646;
    wire N__22645;
    wire N__22644;
    wire N__22643;
    wire N__22642;
    wire N__22641;
    wire N__22640;
    wire N__22639;
    wire N__22638;
    wire N__22637;
    wire N__22636;
    wire N__22635;
    wire N__22634;
    wire N__22633;
    wire N__22632;
    wire N__22631;
    wire N__22630;
    wire N__22629;
    wire N__22628;
    wire N__22627;
    wire N__22626;
    wire N__22625;
    wire N__22624;
    wire N__22623;
    wire N__22622;
    wire N__22621;
    wire N__22620;
    wire N__22619;
    wire N__22618;
    wire N__22617;
    wire N__22616;
    wire N__22615;
    wire N__22614;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22422;
    wire N__22421;
    wire N__22420;
    wire N__22417;
    wire N__22416;
    wire N__22415;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22407;
    wire N__22406;
    wire N__22403;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22379;
    wire N__22378;
    wire N__22373;
    wire N__22370;
    wire N__22365;
    wire N__22360;
    wire N__22355;
    wire N__22352;
    wire N__22339;
    wire N__22336;
    wire N__22335;
    wire N__22334;
    wire N__22333;
    wire N__22332;
    wire N__22331;
    wire N__22328;
    wire N__22327;
    wire N__22326;
    wire N__22325;
    wire N__22324;
    wire N__22323;
    wire N__22320;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22312;
    wire N__22309;
    wire N__22306;
    wire N__22305;
    wire N__22304;
    wire N__22303;
    wire N__22302;
    wire N__22301;
    wire N__22298;
    wire N__22297;
    wire N__22296;
    wire N__22293;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22275;
    wire N__22270;
    wire N__22269;
    wire N__22268;
    wire N__22263;
    wire N__22260;
    wire N__22259;
    wire N__22258;
    wire N__22257;
    wire N__22254;
    wire N__22253;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22231;
    wire N__22226;
    wire N__22221;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22192;
    wire N__22191;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22177;
    wire N__22172;
    wire N__22169;
    wire N__22160;
    wire N__22153;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22135;
    wire N__22130;
    wire N__22125;
    wire N__22120;
    wire N__22115;
    wire N__22102;
    wire N__22101;
    wire N__22100;
    wire N__22097;
    wire N__22096;
    wire N__22095;
    wire N__22094;
    wire N__22093;
    wire N__22092;
    wire N__22091;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22077;
    wire N__22074;
    wire N__22073;
    wire N__22070;
    wire N__22069;
    wire N__22066;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22051;
    wire N__22046;
    wire N__22041;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22014;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21990;
    wire N__21985;
    wire N__21976;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21955;
    wire N__21952;
    wire N__21951;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21947;
    wire N__21944;
    wire N__21943;
    wire N__21942;
    wire N__21941;
    wire N__21938;
    wire N__21933;
    wire N__21930;
    wire N__21929;
    wire N__21928;
    wire N__21927;
    wire N__21924;
    wire N__21923;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21879;
    wire N__21874;
    wire N__21871;
    wire N__21870;
    wire N__21869;
    wire N__21868;
    wire N__21867;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21830;
    wire N__21823;
    wire N__21820;
    wire N__21815;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21792;
    wire N__21791;
    wire N__21790;
    wire N__21789;
    wire N__21788;
    wire N__21787;
    wire N__21784;
    wire N__21783;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21771;
    wire N__21770;
    wire N__21769;
    wire N__21768;
    wire N__21767;
    wire N__21766;
    wire N__21765;
    wire N__21764;
    wire N__21763;
    wire N__21762;
    wire N__21761;
    wire N__21760;
    wire N__21757;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21743;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21716;
    wire N__21715;
    wire N__21714;
    wire N__21707;
    wire N__21702;
    wire N__21699;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21677;
    wire N__21674;
    wire N__21673;
    wire N__21670;
    wire N__21669;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21651;
    wire N__21646;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21628;
    wire N__21625;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21602;
    wire N__21593;
    wire N__21588;
    wire N__21581;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21530;
    wire N__21529;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21515;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21479;
    wire N__21478;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21464;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21444;
    wire N__21441;
    wire N__21440;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21432;
    wire N__21429;
    wire N__21428;
    wire N__21427;
    wire N__21426;
    wire N__21425;
    wire N__21424;
    wire N__21421;
    wire N__21420;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21409;
    wire N__21408;
    wire N__21407;
    wire N__21402;
    wire N__21401;
    wire N__21400;
    wire N__21399;
    wire N__21398;
    wire N__21397;
    wire N__21392;
    wire N__21389;
    wire N__21388;
    wire N__21383;
    wire N__21378;
    wire N__21377;
    wire N__21376;
    wire N__21369;
    wire N__21364;
    wire N__21363;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21351;
    wire N__21344;
    wire N__21341;
    wire N__21336;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21313;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21291;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21277;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21253;
    wire N__21250;
    wire N__21249;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21207;
    wire N__21206;
    wire N__21203;
    wire N__21202;
    wire N__21201;
    wire N__21200;
    wire N__21197;
    wire N__21196;
    wire N__21195;
    wire N__21192;
    wire N__21191;
    wire N__21190;
    wire N__21189;
    wire N__21186;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21175;
    wire N__21174;
    wire N__21173;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21165;
    wire N__21162;
    wire N__21161;
    wire N__21160;
    wire N__21157;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21138;
    wire N__21135;
    wire N__21130;
    wire N__21129;
    wire N__21128;
    wire N__21127;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21109;
    wire N__21104;
    wire N__21095;
    wire N__21092;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21059;
    wire N__21054;
    wire N__21047;
    wire N__21042;
    wire N__21025;
    wire N__21024;
    wire N__21023;
    wire N__21022;
    wire N__21021;
    wire N__21020;
    wire N__21019;
    wire N__21016;
    wire N__21015;
    wire N__21014;
    wire N__21013;
    wire N__21012;
    wire N__21011;
    wire N__21008;
    wire N__21007;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20992;
    wire N__20991;
    wire N__20990;
    wire N__20989;
    wire N__20988;
    wire N__20987;
    wire N__20986;
    wire N__20985;
    wire N__20984;
    wire N__20983;
    wire N__20982;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20964;
    wire N__20961;
    wire N__20956;
    wire N__20953;
    wire N__20948;
    wire N__20945;
    wire N__20940;
    wire N__20937;
    wire N__20932;
    wire N__20931;
    wire N__20930;
    wire N__20929;
    wire N__20928;
    wire N__20927;
    wire N__20920;
    wire N__20913;
    wire N__20912;
    wire N__20911;
    wire N__20910;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20892;
    wire N__20883;
    wire N__20878;
    wire N__20871;
    wire N__20866;
    wire N__20861;
    wire N__20854;
    wire N__20847;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20814;
    wire N__20811;
    wire N__20810;
    wire N__20809;
    wire N__20808;
    wire N__20807;
    wire N__20806;
    wire N__20805;
    wire N__20804;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20792;
    wire N__20791;
    wire N__20788;
    wire N__20787;
    wire N__20786;
    wire N__20785;
    wire N__20784;
    wire N__20781;
    wire N__20776;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20758;
    wire N__20757;
    wire N__20754;
    wire N__20753;
    wire N__20752;
    wire N__20749;
    wire N__20742;
    wire N__20737;
    wire N__20734;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20719;
    wire N__20718;
    wire N__20717;
    wire N__20714;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20697;
    wire N__20692;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20671;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20631;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20611;
    wire N__20608;
    wire N__20603;
    wire N__20600;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20577;
    wire N__20576;
    wire N__20575;
    wire N__20574;
    wire N__20573;
    wire N__20572;
    wire N__20571;
    wire N__20570;
    wire N__20569;
    wire N__20566;
    wire N__20565;
    wire N__20564;
    wire N__20563;
    wire N__20562;
    wire N__20557;
    wire N__20556;
    wire N__20555;
    wire N__20554;
    wire N__20551;
    wire N__20544;
    wire N__20541;
    wire N__20540;
    wire N__20539;
    wire N__20538;
    wire N__20537;
    wire N__20532;
    wire N__20531;
    wire N__20530;
    wire N__20527;
    wire N__20522;
    wire N__20521;
    wire N__20516;
    wire N__20513;
    wire N__20512;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20492;
    wire N__20489;
    wire N__20488;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20463;
    wire N__20462;
    wire N__20459;
    wire N__20458;
    wire N__20455;
    wire N__20454;
    wire N__20451;
    wire N__20444;
    wire N__20443;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20404;
    wire N__20401;
    wire N__20396;
    wire N__20391;
    wire N__20382;
    wire N__20365;
    wire N__20364;
    wire N__20363;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20349;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20320;
    wire N__20317;
    wire N__20312;
    wire N__20309;
    wire N__20308;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20284;
    wire N__20283;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20272;
    wire N__20271;
    wire N__20270;
    wire N__20269;
    wire N__20268;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20257;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20230;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20209;
    wire N__20206;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20188;
    wire N__20185;
    wire N__20184;
    wire N__20179;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20164;
    wire N__20163;
    wire N__20156;
    wire N__20155;
    wire N__20152;
    wire N__20147;
    wire N__20144;
    wire N__20137;
    wire N__20132;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20116;
    wire N__20111;
    wire N__20098;
    wire N__20097;
    wire N__20096;
    wire N__20095;
    wire N__20094;
    wire N__20093;
    wire N__20092;
    wire N__20091;
    wire N__20090;
    wire N__20089;
    wire N__20088;
    wire N__20085;
    wire N__20084;
    wire N__20083;
    wire N__20082;
    wire N__20081;
    wire N__20080;
    wire N__20079;
    wire N__20078;
    wire N__20077;
    wire N__20076;
    wire N__20075;
    wire N__20072;
    wire N__20071;
    wire N__20070;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20062;
    wire N__20061;
    wire N__20060;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20052;
    wire N__20051;
    wire N__20050;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20028;
    wire N__20021;
    wire N__20020;
    wire N__20019;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20002;
    wire N__19999;
    wire N__19998;
    wire N__19997;
    wire N__19996;
    wire N__19993;
    wire N__19992;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19978;
    wire N__19973;
    wire N__19972;
    wire N__19971;
    wire N__19970;
    wire N__19969;
    wire N__19968;
    wire N__19967;
    wire N__19966;
    wire N__19965;
    wire N__19964;
    wire N__19963;
    wire N__19962;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19944;
    wire N__19941;
    wire N__19936;
    wire N__19931;
    wire N__19928;
    wire N__19923;
    wire N__19918;
    wire N__19917;
    wire N__19916;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19904;
    wire N__19899;
    wire N__19894;
    wire N__19889;
    wire N__19886;
    wire N__19881;
    wire N__19880;
    wire N__19879;
    wire N__19878;
    wire N__19877;
    wire N__19876;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19857;
    wire N__19850;
    wire N__19847;
    wire N__19836;
    wire N__19835;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19821;
    wire N__19814;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19796;
    wire N__19793;
    wire N__19788;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19762;
    wire N__19757;
    wire N__19752;
    wire N__19743;
    wire N__19736;
    wire N__19717;
    wire N__19716;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19704;
    wire N__19703;
    wire N__19700;
    wire N__19699;
    wire N__19698;
    wire N__19697;
    wire N__19696;
    wire N__19695;
    wire N__19692;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19680;
    wire N__19679;
    wire N__19678;
    wire N__19675;
    wire N__19670;
    wire N__19667;
    wire N__19666;
    wire N__19663;
    wire N__19662;
    wire N__19659;
    wire N__19658;
    wire N__19655;
    wire N__19654;
    wire N__19651;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19632;
    wire N__19629;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19605;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19579;
    wire N__19574;
    wire N__19561;
    wire N__19560;
    wire N__19557;
    wire N__19556;
    wire N__19555;
    wire N__19554;
    wire N__19553;
    wire N__19552;
    wire N__19551;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19539;
    wire N__19538;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19530;
    wire N__19525;
    wire N__19522;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19487;
    wire N__19486;
    wire N__19485;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19450;
    wire N__19447;
    wire N__19440;
    wire N__19429;
    wire N__19426;
    wire N__19425;
    wire N__19422;
    wire N__19419;
    wire N__19416;
    wire N__19413;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19380;
    wire N__19379;
    wire N__19372;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19360;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19348;
    wire N__19345;
    wire N__19344;
    wire N__19343;
    wire N__19342;
    wire N__19335;
    wire N__19332;
    wire N__19327;
    wire N__19324;
    wire N__19323;
    wire N__19320;
    wire N__19319;
    wire N__19316;
    wire N__19315;
    wire N__19314;
    wire N__19311;
    wire N__19310;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19293;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19254;
    wire N__19243;
    wire N__19240;
    wire N__19239;
    wire N__19238;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19220;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19212;
    wire N__19211;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19199;
    wire N__19194;
    wire N__19191;
    wire N__19180;
    wire N__19177;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19167;
    wire N__19166;
    wire N__19165;
    wire N__19164;
    wire N__19163;
    wire N__19162;
    wire N__19161;
    wire N__19158;
    wire N__19157;
    wire N__19156;
    wire N__19155;
    wire N__19152;
    wire N__19151;
    wire N__19150;
    wire N__19149;
    wire N__19148;
    wire N__19147;
    wire N__19144;
    wire N__19139;
    wire N__19134;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19118;
    wire N__19113;
    wire N__19110;
    wire N__19109;
    wire N__19108;
    wire N__19107;
    wire N__19102;
    wire N__19101;
    wire N__19098;
    wire N__19097;
    wire N__19096;
    wire N__19091;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19041;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19027;
    wire N__19022;
    wire N__19017;
    wire N__19010;
    wire N__19003;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18954;
    wire N__18953;
    wire N__18952;
    wire N__18951;
    wire N__18948;
    wire N__18947;
    wire N__18946;
    wire N__18943;
    wire N__18940;
    wire N__18939;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18922;
    wire N__18919;
    wire N__18918;
    wire N__18915;
    wire N__18914;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18869;
    wire N__18864;
    wire N__18859;
    wire N__18858;
    wire N__18855;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18833;
    wire N__18830;
    wire N__18823;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18783;
    wire N__18782;
    wire N__18781;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18773;
    wire N__18772;
    wire N__18771;
    wire N__18766;
    wire N__18765;
    wire N__18764;
    wire N__18763;
    wire N__18760;
    wire N__18755;
    wire N__18752;
    wire N__18751;
    wire N__18750;
    wire N__18749;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18731;
    wire N__18730;
    wire N__18729;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18721;
    wire N__18720;
    wire N__18719;
    wire N__18716;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18684;
    wire N__18679;
    wire N__18672;
    wire N__18667;
    wire N__18658;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18627;
    wire N__18626;
    wire N__18625;
    wire N__18624;
    wire N__18623;
    wire N__18622;
    wire N__18621;
    wire N__18620;
    wire N__18617;
    wire N__18616;
    wire N__18613;
    wire N__18612;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18602;
    wire N__18601;
    wire N__18600;
    wire N__18599;
    wire N__18592;
    wire N__18591;
    wire N__18590;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18580;
    wire N__18573;
    wire N__18572;
    wire N__18571;
    wire N__18566;
    wire N__18563;
    wire N__18562;
    wire N__18559;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18532;
    wire N__18529;
    wire N__18524;
    wire N__18519;
    wire N__18512;
    wire N__18507;
    wire N__18504;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18443;
    wire N__18442;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18426;
    wire N__18423;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18340;
    wire N__18337;
    wire N__18336;
    wire N__18333;
    wire N__18332;
    wire N__18331;
    wire N__18328;
    wire N__18327;
    wire N__18326;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18316;
    wire N__18315;
    wire N__18310;
    wire N__18309;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18247;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18236;
    wire N__18231;
    wire N__18228;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18199;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18165;
    wire N__18164;
    wire N__18157;
    wire N__18156;
    wire N__18155;
    wire N__18152;
    wire N__18147;
    wire N__18142;
    wire N__18141;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18091;
    wire N__18088;
    wire N__18087;
    wire N__18086;
    wire N__18085;
    wire N__18084;
    wire N__18083;
    wire N__18082;
    wire N__18081;
    wire N__18080;
    wire N__18079;
    wire N__18078;
    wire N__18077;
    wire N__18076;
    wire N__18075;
    wire N__18074;
    wire N__18073;
    wire N__18072;
    wire N__18071;
    wire N__18070;
    wire N__18069;
    wire N__18068;
    wire N__18067;
    wire N__18066;
    wire N__18065;
    wire N__18064;
    wire N__18063;
    wire N__18062;
    wire N__18061;
    wire N__18060;
    wire N__18059;
    wire N__18058;
    wire N__18057;
    wire N__18056;
    wire N__18055;
    wire N__18054;
    wire N__18053;
    wire N__18052;
    wire N__18051;
    wire N__18050;
    wire N__18049;
    wire N__18048;
    wire N__18047;
    wire N__18046;
    wire N__18045;
    wire N__18044;
    wire N__18043;
    wire N__18042;
    wire N__18041;
    wire N__18040;
    wire N__18039;
    wire N__18038;
    wire N__18035;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17925;
    wire N__17922;
    wire N__17919;
    wire N__17916;
    wire N__17913;
    wire N__17908;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17898;
    wire N__17897;
    wire N__17894;
    wire N__17889;
    wire N__17888;
    wire N__17883;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17863;
    wire N__17860;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17848;
    wire N__17845;
    wire N__17842;
    wire N__17841;
    wire N__17840;
    wire N__17839;
    wire N__17838;
    wire N__17833;
    wire N__17832;
    wire N__17831;
    wire N__17830;
    wire N__17829;
    wire N__17826;
    wire N__17821;
    wire N__17818;
    wire N__17811;
    wire N__17810;
    wire N__17809;
    wire N__17808;
    wire N__17807;
    wire N__17802;
    wire N__17799;
    wire N__17794;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17773;
    wire N__17768;
    wire N__17765;
    wire N__17762;
    wire N__17757;
    wire N__17752;
    wire N__17749;
    wire N__17746;
    wire N__17743;
    wire N__17740;
    wire N__17737;
    wire N__17734;
    wire N__17731;
    wire N__17730;
    wire N__17727;
    wire N__17724;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17709;
    wire N__17708;
    wire N__17705;
    wire N__17700;
    wire N__17695;
    wire N__17692;
    wire N__17691;
    wire N__17688;
    wire N__17687;
    wire N__17686;
    wire N__17685;
    wire N__17682;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17655;
    wire N__17652;
    wire N__17645;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17625;
    wire N__17624;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17616;
    wire N__17615;
    wire N__17612;
    wire N__17611;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17577;
    wire N__17576;
    wire N__17575;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17554;
    wire N__17551;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17524;
    wire N__17521;
    wire N__17520;
    wire N__17517;
    wire N__17514;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17502;
    wire N__17501;
    wire N__17500;
    wire N__17499;
    wire N__17498;
    wire N__17497;
    wire N__17496;
    wire N__17495;
    wire N__17494;
    wire N__17491;
    wire N__17490;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17482;
    wire N__17477;
    wire N__17476;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17446;
    wire N__17443;
    wire N__17442;
    wire N__17441;
    wire N__17440;
    wire N__17437;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17417;
    wire N__17412;
    wire N__17409;
    wire N__17406;
    wire N__17401;
    wire N__17398;
    wire N__17393;
    wire N__17388;
    wire N__17383;
    wire N__17368;
    wire N__17367;
    wire N__17364;
    wire N__17363;
    wire N__17360;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17336;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17310;
    wire N__17299;
    wire N__17296;
    wire N__17293;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17217;
    wire N__17216;
    wire N__17215;
    wire N__17212;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17182;
    wire N__17179;
    wire N__17178;
    wire N__17175;
    wire N__17174;
    wire N__17171;
    wire N__17170;
    wire N__17167;
    wire N__17160;
    wire N__17155;
    wire N__17154;
    wire N__17151;
    wire N__17150;
    wire N__17149;
    wire N__17148;
    wire N__17145;
    wire N__17136;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17112;
    wire N__17111;
    wire N__17110;
    wire N__17107;
    wire N__17100;
    wire N__17095;
    wire N__17092;
    wire N__17091;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17076;
    wire N__17075;
    wire N__17074;
    wire N__17073;
    wire N__17072;
    wire N__17067;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17049;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17031;
    wire N__17028;
    wire N__17023;
    wire N__17022;
    wire N__17021;
    wire N__17020;
    wire N__17019;
    wire N__17016;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__16999;
    wire N__16994;
    wire N__16989;
    wire N__16972;
    wire N__16971;
    wire N__16970;
    wire N__16967;
    wire N__16966;
    wire N__16965;
    wire N__16964;
    wire N__16961;
    wire N__16960;
    wire N__16959;
    wire N__16958;
    wire N__16957;
    wire N__16956;
    wire N__16955;
    wire N__16954;
    wire N__16951;
    wire N__16946;
    wire N__16945;
    wire N__16944;
    wire N__16943;
    wire N__16942;
    wire N__16941;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16921;
    wire N__16918;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16906;
    wire N__16901;
    wire N__16900;
    wire N__16899;
    wire N__16896;
    wire N__16891;
    wire N__16890;
    wire N__16887;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16879;
    wire N__16878;
    wire N__16877;
    wire N__16874;
    wire N__16867;
    wire N__16864;
    wire N__16855;
    wire N__16854;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16846;
    wire N__16843;
    wire N__16840;
    wire N__16833;
    wire N__16828;
    wire N__16825;
    wire N__16820;
    wire N__16815;
    wire N__16810;
    wire N__16801;
    wire N__16798;
    wire N__16791;
    wire N__16774;
    wire N__16771;
    wire N__16768;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16758;
    wire N__16757;
    wire N__16756;
    wire N__16755;
    wire N__16754;
    wire N__16753;
    wire N__16752;
    wire N__16735;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16708;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16696;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16678;
    wire N__16675;
    wire N__16672;
    wire N__16669;
    wire N__16668;
    wire N__16667;
    wire N__16664;
    wire N__16659;
    wire N__16656;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16642;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16623;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16605;
    wire N__16604;
    wire N__16603;
    wire N__16600;
    wire N__16593;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16581;
    wire N__16578;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16561;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16550;
    wire N__16549;
    wire N__16548;
    wire N__16547;
    wire N__16546;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16527;
    wire N__16520;
    wire N__16513;
    wire N__16510;
    wire N__16509;
    wire N__16506;
    wire N__16505;
    wire N__16504;
    wire N__16501;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16490;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16463;
    wire N__16450;
    wire N__16447;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16437;
    wire N__16434;
    wire N__16433;
    wire N__16432;
    wire N__16427;
    wire N__16422;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16405;
    wire N__16402;
    wire N__16399;
    wire N__16396;
    wire N__16393;
    wire N__16390;
    wire N__16387;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16371;
    wire N__16368;
    wire N__16367;
    wire N__16364;
    wire N__16359;
    wire N__16358;
    wire N__16355;
    wire N__16354;
    wire N__16353;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16343;
    wire N__16342;
    wire N__16341;
    wire N__16338;
    wire N__16333;
    wire N__16330;
    wire N__16327;
    wire N__16324;
    wire N__16319;
    wire N__16306;
    wire N__16305;
    wire N__16304;
    wire N__16301;
    wire N__16298;
    wire N__16297;
    wire N__16294;
    wire N__16293;
    wire N__16292;
    wire N__16291;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16256;
    wire N__16251;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16230;
    wire N__16227;
    wire N__16224;
    wire N__16221;
    wire N__16218;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16185;
    wire N__16184;
    wire N__16181;
    wire N__16176;
    wire N__16171;
    wire N__16170;
    wire N__16169;
    wire N__16168;
    wire N__16167;
    wire N__16166;
    wire N__16165;
    wire N__16164;
    wire N__16163;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16155;
    wire N__16150;
    wire N__16147;
    wire N__16146;
    wire N__16143;
    wire N__16142;
    wire N__16137;
    wire N__16136;
    wire N__16133;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16104;
    wire N__16101;
    wire N__16096;
    wire N__16089;
    wire N__16076;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16021;
    wire N__16018;
    wire N__16015;
    wire N__16012;
    wire N__16009;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15985;
    wire N__15984;
    wire N__15981;
    wire N__15978;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15945;
    wire N__15944;
    wire N__15943;
    wire N__15936;
    wire N__15933;
    wire N__15928;
    wire N__15925;
    wire N__15924;
    wire N__15923;
    wire N__15922;
    wire N__15915;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15905;
    wire N__15898;
    wire N__15897;
    wire N__15896;
    wire N__15895;
    wire N__15892;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15878;
    wire N__15875;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15858;
    wire N__15857;
    wire N__15856;
    wire N__15853;
    wire N__15848;
    wire N__15845;
    wire N__15838;
    wire N__15835;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15820;
    wire N__15819;
    wire N__15818;
    wire N__15813;
    wire N__15810;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15793;
    wire N__15790;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15782;
    wire N__15777;
    wire N__15776;
    wire N__15773;
    wire N__15772;
    wire N__15771;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15759;
    wire N__15758;
    wire N__15755;
    wire N__15754;
    wire N__15753;
    wire N__15752;
    wire N__15747;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15728;
    wire N__15723;
    wire N__15720;
    wire N__15717;
    wire N__15706;
    wire N__15705;
    wire N__15704;
    wire N__15703;
    wire N__15702;
    wire N__15697;
    wire N__15696;
    wire N__15695;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15687;
    wire N__15686;
    wire N__15683;
    wire N__15682;
    wire N__15681;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15666;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15652;
    wire N__15651;
    wire N__15650;
    wire N__15647;
    wire N__15642;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15607;
    wire N__15602;
    wire N__15593;
    wire N__15588;
    wire N__15581;
    wire N__15568;
    wire N__15567;
    wire N__15562;
    wire N__15561;
    wire N__15560;
    wire N__15559;
    wire N__15558;
    wire N__15557;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15541;
    wire N__15538;
    wire N__15529;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15514;
    wire N__15511;
    wire N__15510;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15499;
    wire N__15498;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15490;
    wire N__15489;
    wire N__15482;
    wire N__15479;
    wire N__15474;
    wire N__15469;
    wire N__15464;
    wire N__15461;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15447;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15433;
    wire N__15432;
    wire N__15431;
    wire N__15430;
    wire N__15429;
    wire N__15426;
    wire N__15417;
    wire N__15412;
    wire N__15411;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15399;
    wire N__15396;
    wire N__15391;
    wire N__15390;
    wire N__15387;
    wire N__15386;
    wire N__15385;
    wire N__15384;
    wire N__15383;
    wire N__15380;
    wire N__15369;
    wire N__15366;
    wire N__15365;
    wire N__15364;
    wire N__15361;
    wire N__15358;
    wire N__15353;
    wire N__15350;
    wire N__15343;
    wire N__15340;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15325;
    wire N__15324;
    wire N__15323;
    wire N__15322;
    wire N__15321;
    wire N__15318;
    wire N__15317;
    wire N__15316;
    wire N__15313;
    wire N__15306;
    wire N__15303;
    wire N__15298;
    wire N__15291;
    wire N__15286;
    wire N__15283;
    wire N__15282;
    wire N__15281;
    wire N__15280;
    wire N__15279;
    wire N__15278;
    wire N__15277;
    wire N__15276;
    wire N__15275;
    wire N__15274;
    wire N__15273;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15265;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15252;
    wire N__15251;
    wire N__15250;
    wire N__15249;
    wire N__15248;
    wire N__15247;
    wire N__15244;
    wire N__15241;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15233;
    wire N__15232;
    wire N__15231;
    wire N__15230;
    wire N__15229;
    wire N__15228;
    wire N__15225;
    wire N__15224;
    wire N__15223;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15184;
    wire N__15183;
    wire N__15182;
    wire N__15175;
    wire N__15158;
    wire N__15151;
    wire N__15148;
    wire N__15143;
    wire N__15140;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15118;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15104;
    wire N__15101;
    wire N__15082;
    wire N__15081;
    wire N__15078;
    wire N__15077;
    wire N__15076;
    wire N__15075;
    wire N__15072;
    wire N__15069;
    wire N__15066;
    wire N__15061;
    wire N__15052;
    wire N__15049;
    wire N__15048;
    wire N__15045;
    wire N__15042;
    wire N__15039;
    wire N__15034;
    wire N__15031;
    wire N__15030;
    wire N__15027;
    wire N__15024;
    wire N__15021;
    wire N__15018;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__15001;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14985;
    wire N__14984;
    wire N__14983;
    wire N__14982;
    wire N__14981;
    wire N__14980;
    wire N__14973;
    wire N__14970;
    wire N__14967;
    wire N__14964;
    wire N__14961;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14943;
    wire N__14940;
    wire N__14937;
    wire N__14934;
    wire N__14929;
    wire N__14928;
    wire N__14925;
    wire N__14922;
    wire N__14919;
    wire N__14914;
    wire N__14911;
    wire N__14910;
    wire N__14909;
    wire N__14908;
    wire N__14905;
    wire N__14898;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14872;
    wire N__14869;
    wire N__14868;
    wire N__14867;
    wire N__14866;
    wire N__14863;
    wire N__14856;
    wire N__14855;
    wire N__14854;
    wire N__14849;
    wire N__14846;
    wire N__14845;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14830;
    wire N__14827;
    wire N__14818;
    wire N__14815;
    wire N__14814;
    wire N__14809;
    wire N__14806;
    wire N__14805;
    wire N__14802;
    wire N__14799;
    wire N__14794;
    wire N__14793;
    wire N__14792;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14762;
    wire N__14757;
    wire N__14752;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14737;
    wire N__14734;
    wire N__14731;
    wire N__14728;
    wire N__14727;
    wire N__14724;
    wire N__14721;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14680;
    wire N__14677;
    wire N__14676;
    wire N__14673;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14622;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14602;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14538;
    wire N__14537;
    wire N__14536;
    wire N__14533;
    wire N__14526;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14475;
    wire N__14474;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14464;
    wire N__14461;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14442;
    wire N__14439;
    wire N__14434;
    wire N__14433;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14421;
    wire N__14418;
    wire N__14415;
    wire N__14410;
    wire N__14407;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14346;
    wire N__14343;
    wire N__14340;
    wire N__14335;
    wire N__14332;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14310;
    wire N__14305;
    wire N__14302;
    wire N__14301;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14242;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14199;
    wire N__14198;
    wire N__14195;
    wire N__14194;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14169;
    wire N__14166;
    wire N__14163;
    wire N__14160;
    wire N__14155;
    wire N__14154;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14146;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14124;
    wire N__14119;
    wire N__14118;
    wire N__14117;
    wire N__14114;
    wire N__14109;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14087;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14069;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14040;
    wire N__14037;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14023;
    wire N__14020;
    wire N__14019;
    wire N__14014;
    wire N__14013;
    wire N__14010;
    wire N__14007;
    wire N__14002;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13989;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13966;
    wire N__13965;
    wire N__13964;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13923;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13911;
    wire N__13908;
    wire N__13905;
    wire N__13900;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13885;
    wire N__13884;
    wire N__13879;
    wire N__13876;
    wire N__13873;
    wire N__13870;
    wire N__13869;
    wire N__13866;
    wire N__13863;
    wire N__13860;
    wire N__13855;
    wire N__13852;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13837;
    wire N__13836;
    wire N__13835;
    wire N__13834;
    wire N__13831;
    wire N__13828;
    wire N__13823;
    wire N__13816;
    wire N__13815;
    wire N__13812;
    wire N__13809;
    wire N__13806;
    wire N__13803;
    wire N__13800;
    wire N__13795;
    wire N__13792;
    wire N__13791;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13779;
    wire N__13776;
    wire N__13771;
    wire N__13770;
    wire N__13769;
    wire N__13768;
    wire N__13767;
    wire N__13764;
    wire N__13759;
    wire N__13754;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13726;
    wire N__13725;
    wire N__13724;
    wire N__13723;
    wire N__13722;
    wire N__13719;
    wire N__13714;
    wire N__13711;
    wire N__13708;
    wire N__13699;
    wire N__13696;
    wire N__13695;
    wire N__13692;
    wire N__13689;
    wire N__13686;
    wire N__13681;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13669;
    wire N__13666;
    wire N__13665;
    wire N__13662;
    wire N__13659;
    wire N__13654;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13644;
    wire N__13639;
    wire N__13638;
    wire N__13637;
    wire N__13636;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13621;
    wire N__13618;
    wire N__13609;
    wire N__13606;
    wire N__13603;
    wire N__13602;
    wire N__13599;
    wire N__13596;
    wire N__13593;
    wire N__13588;
    wire N__13585;
    wire N__13584;
    wire N__13583;
    wire N__13580;
    wire N__13575;
    wire N__13572;
    wire N__13567;
    wire N__13564;
    wire N__13561;
    wire N__13558;
    wire N__13555;
    wire N__13552;
    wire N__13549;
    wire N__13546;
    wire N__13543;
    wire N__13540;
    wire N__13537;
    wire N__13534;
    wire N__13531;
    wire N__13528;
    wire N__13525;
    wire N__13522;
    wire N__13519;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13495;
    wire N__13492;
    wire N__13489;
    wire N__13486;
    wire N__13483;
    wire N__13482;
    wire N__13477;
    wire N__13474;
    wire N__13473;
    wire N__13470;
    wire N__13469;
    wire N__13468;
    wire N__13465;
    wire N__13464;
    wire N__13461;
    wire N__13456;
    wire N__13453;
    wire N__13450;
    wire N__13447;
    wire N__13438;
    wire N__13437;
    wire N__13434;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13413;
    wire N__13412;
    wire N__13411;
    wire N__13410;
    wire N__13409;
    wire N__13408;
    wire N__13407;
    wire N__13406;
    wire N__13401;
    wire N__13396;
    wire N__13385;
    wire N__13378;
    wire N__13377;
    wire N__13376;
    wire N__13375;
    wire N__13374;
    wire N__13373;
    wire N__13370;
    wire N__13365;
    wire N__13358;
    wire N__13357;
    wire N__13354;
    wire N__13351;
    wire N__13350;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13338;
    wire N__13333;
    wire N__13324;
    wire N__13323;
    wire N__13322;
    wire N__13319;
    wire N__13318;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13305;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13291;
    wire N__13288;
    wire N__13279;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13267;
    wire N__13264;
    wire N__13261;
    wire N__13258;
    wire N__13255;
    wire N__13252;
    wire N__13251;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13219;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13207;
    wire N__13204;
    wire N__13201;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13189;
    wire N__13186;
    wire N__13183;
    wire N__13182;
    wire N__13181;
    wire N__13174;
    wire N__13171;
    wire N__13170;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13156;
    wire N__13153;
    wire N__13150;
    wire N__13147;
    wire N__13146;
    wire N__13143;
    wire N__13140;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13126;
    wire N__13123;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13110;
    wire N__13105;
    wire N__13102;
    wire N__13099;
    wire N__13096;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13086;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13069;
    wire N__13066;
    wire N__13063;
    wire N__13060;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13048;
    wire N__13045;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13035;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13017;
    wire N__13016;
    wire N__13013;
    wire N__13010;
    wire N__13007;
    wire N__13000;
    wire N__12997;
    wire N__12994;
    wire N__12991;
    wire N__12988;
    wire N__12985;
    wire N__12982;
    wire N__12979;
    wire N__12976;
    wire N__12973;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12961;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12951;
    wire N__12946;
    wire N__12945;
    wire N__12942;
    wire N__12939;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12927;
    wire N__12922;
    wire N__12919;
    wire N__12916;
    wire N__12913;
    wire N__12910;
    wire N__12907;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12886;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12865;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12841;
    wire N__12838;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12823;
    wire N__12820;
    wire N__12819;
    wire N__12816;
    wire N__12813;
    wire N__12810;
    wire N__12807;
    wire N__12802;
    wire N__12801;
    wire N__12800;
    wire N__12799;
    wire N__12798;
    wire N__12797;
    wire N__12796;
    wire N__12795;
    wire N__12794;
    wire N__12793;
    wire N__12792;
    wire N__12791;
    wire N__12790;
    wire N__12789;
    wire N__12788;
    wire N__12787;
    wire N__12786;
    wire N__12769;
    wire N__12752;
    wire N__12751;
    wire N__12750;
    wire N__12749;
    wire N__12748;
    wire N__12747;
    wire N__12746;
    wire N__12745;
    wire N__12744;
    wire N__12743;
    wire N__12742;
    wire N__12741;
    wire N__12740;
    wire N__12739;
    wire N__12738;
    wire N__12737;
    wire N__12736;
    wire N__12733;
    wire N__12728;
    wire N__12713;
    wire N__12710;
    wire N__12693;
    wire N__12688;
    wire N__12683;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12655;
    wire N__12654;
    wire N__12651;
    wire N__12648;
    wire N__12645;
    wire N__12640;
    wire N__12637;
    wire N__12634;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12598;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12582;
    wire N__12577;
    wire N__12574;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12559;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12549;
    wire N__12544;
    wire N__12541;
    wire N__12540;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12526;
    wire N__12523;
    wire N__12522;
    wire N__12519;
    wire N__12516;
    wire N__12513;
    wire N__12508;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12500;
    wire N__12497;
    wire N__12492;
    wire N__12489;
    wire N__12484;
    wire N__12483;
    wire N__12480;
    wire N__12477;
    wire N__12474;
    wire N__12469;
    wire N__12468;
    wire N__12467;
    wire N__12466;
    wire N__12457;
    wire N__12454;
    wire N__12451;
    wire N__12450;
    wire N__12447;
    wire N__12444;
    wire N__12439;
    wire N__12436;
    wire N__12435;
    wire N__12434;
    wire N__12431;
    wire N__12430;
    wire N__12427;
    wire N__12426;
    wire N__12425;
    wire N__12424;
    wire N__12423;
    wire N__12420;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12405;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12379;
    wire N__12376;
    wire N__12373;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12361;
    wire N__12358;
    wire N__12357;
    wire N__12356;
    wire N__12353;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12337;
    wire N__12334;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12313;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12305;
    wire N__12304;
    wire N__12299;
    wire N__12294;
    wire N__12291;
    wire N__12286;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12276;
    wire N__12271;
    wire N__12268;
    wire N__12267;
    wire N__12264;
    wire N__12263;
    wire N__12260;
    wire N__12259;
    wire N__12258;
    wire N__12255;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12237;
    wire N__12232;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12219;
    wire N__12216;
    wire N__12213;
    wire N__12208;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12198;
    wire N__12195;
    wire N__12192;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12180;
    wire N__12179;
    wire N__12178;
    wire N__12177;
    wire N__12176;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12159;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12132;
    wire N__12127;
    wire N__12124;
    wire N__12115;
    wire N__12112;
    wire N__12109;
    wire N__12106;
    wire N__12105;
    wire N__12104;
    wire N__12103;
    wire N__12100;
    wire N__12097;
    wire N__12096;
    wire N__12095;
    wire N__12094;
    wire N__12093;
    wire N__12090;
    wire N__12087;
    wire N__12086;
    wire N__12081;
    wire N__12078;
    wire N__12071;
    wire N__12064;
    wire N__12059;
    wire N__12052;
    wire N__12051;
    wire N__12050;
    wire N__12049;
    wire N__12048;
    wire N__12047;
    wire N__12044;
    wire N__12043;
    wire N__12042;
    wire N__12041;
    wire N__12040;
    wire N__12039;
    wire N__12038;
    wire N__12037;
    wire N__12036;
    wire N__12035;
    wire N__12030;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12012;
    wire N__12009;
    wire N__12002;
    wire N__11997;
    wire N__11994;
    wire N__11989;
    wire N__11986;
    wire N__11981;
    wire N__11968;
    wire N__11965;
    wire N__11964;
    wire N__11961;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11940;
    wire N__11935;
    wire N__11934;
    wire N__11933;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11925;
    wire N__11924;
    wire N__11923;
    wire N__11922;
    wire N__11921;
    wire N__11914;
    wire N__11911;
    wire N__11904;
    wire N__11899;
    wire N__11898;
    wire N__11897;
    wire N__11894;
    wire N__11887;
    wire N__11882;
    wire N__11877;
    wire N__11872;
    wire N__11869;
    wire N__11866;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11851;
    wire N__11848;
    wire N__11847;
    wire N__11844;
    wire N__11839;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11829;
    wire N__11824;
    wire N__11823;
    wire N__11820;
    wire N__11819;
    wire N__11816;
    wire N__11813;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11797;
    wire N__11796;
    wire N__11793;
    wire N__11790;
    wire N__11787;
    wire N__11782;
    wire N__11779;
    wire N__11778;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11758;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11743;
    wire N__11742;
    wire N__11741;
    wire N__11738;
    wire N__11733;
    wire N__11730;
    wire N__11725;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11689;
    wire N__11686;
    wire N__11683;
    wire N__11680;
    wire N__11679;
    wire N__11678;
    wire N__11675;
    wire N__11674;
    wire N__11669;
    wire N__11666;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11619;
    wire N__11616;
    wire N__11613;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11592;
    wire N__11587;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11562;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11523;
    wire N__11520;
    wire N__11519;
    wire N__11518;
    wire N__11517;
    wire N__11514;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11496;
    wire N__11485;
    wire N__11484;
    wire N__11481;
    wire N__11478;
    wire N__11473;
    wire N__11470;
    wire N__11469;
    wire N__11468;
    wire N__11467;
    wire N__11464;
    wire N__11463;
    wire N__11462;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11452;
    wire N__11449;
    wire N__11444;
    wire N__11443;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11433;
    wire N__11432;
    wire N__11429;
    wire N__11424;
    wire N__11419;
    wire N__11416;
    wire N__11411;
    wire N__11408;
    wire N__11395;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11387;
    wire N__11386;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11375;
    wire N__11374;
    wire N__11371;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11359;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11340;
    wire N__11335;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11319;
    wire N__11316;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11302;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11294;
    wire N__11293;
    wire N__11288;
    wire N__11283;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11268;
    wire N__11267;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11262;
    wire N__11257;
    wire N__11246;
    wire N__11243;
    wire N__11242;
    wire N__11241;
    wire N__11238;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11226;
    wire N__11225;
    wire N__11218;
    wire N__11215;
    wire N__11210;
    wire N__11207;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11184;
    wire N__11183;
    wire N__11180;
    wire N__11175;
    wire N__11170;
    wire N__11169;
    wire N__11164;
    wire N__11161;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11149;
    wire N__11148;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11131;
    wire N__11128;
    wire N__11125;
    wire N__11122;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11107;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11092;
    wire N__11091;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11063;
    wire N__11058;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11044;
    wire N__11041;
    wire N__11040;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11017;
    wire N__11014;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10996;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10981;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10969;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10959;
    wire N__10954;
    wire N__10951;
    wire N__10950;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10932;
    wire N__10927;
    wire N__10926;
    wire N__10923;
    wire N__10920;
    wire N__10915;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10900;
    wire N__10899;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10885;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10875;
    wire N__10870;
    wire N__10869;
    wire N__10866;
    wire N__10863;
    wire N__10860;
    wire N__10857;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10825;
    wire N__10824;
    wire N__10821;
    wire N__10818;
    wire N__10813;
    wire N__10812;
    wire N__10809;
    wire N__10806;
    wire N__10803;
    wire N__10798;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10768;
    wire N__10767;
    wire N__10764;
    wire N__10761;
    wire N__10758;
    wire N__10753;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10738;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10726;
    wire N__10725;
    wire N__10722;
    wire N__10719;
    wire N__10714;
    wire N__10711;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10698;
    wire N__10695;
    wire N__10690;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10678;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10666;
    wire N__10665;
    wire N__10660;
    wire N__10657;
    wire N__10656;
    wire N__10653;
    wire N__10652;
    wire N__10651;
    wire N__10650;
    wire N__10649;
    wire N__10648;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10636;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10609;
    wire N__10608;
    wire N__10605;
    wire N__10604;
    wire N__10603;
    wire N__10600;
    wire N__10599;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10591;
    wire N__10590;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10578;
    wire N__10573;
    wire N__10570;
    wire N__10565;
    wire N__10552;
    wire N__10551;
    wire N__10550;
    wire N__10549;
    wire N__10548;
    wire N__10547;
    wire N__10546;
    wire N__10541;
    wire N__10536;
    wire N__10535;
    wire N__10534;
    wire N__10531;
    wire N__10528;
    wire N__10525;
    wire N__10522;
    wire N__10519;
    wire N__10516;
    wire N__10511;
    wire N__10498;
    wire N__10497;
    wire N__10496;
    wire N__10495;
    wire N__10494;
    wire N__10491;
    wire N__10490;
    wire N__10487;
    wire N__10486;
    wire N__10481;
    wire N__10478;
    wire N__10477;
    wire N__10474;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10460;
    wire N__10457;
    wire N__10444;
    wire N__10441;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10420;
    wire N__10419;
    wire N__10416;
    wire N__10413;
    wire N__10408;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10377;
    wire N__10374;
    wire N__10373;
    wire N__10368;
    wire N__10367;
    wire N__10366;
    wire N__10365;
    wire N__10364;
    wire N__10361;
    wire N__10360;
    wire N__10359;
    wire N__10358;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10346;
    wire N__10343;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10321;
    wire N__10314;
    wire N__10309;
    wire N__10308;
    wire N__10307;
    wire N__10306;
    wire N__10305;
    wire N__10296;
    wire N__10293;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10278;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10266;
    wire N__10263;
    wire N__10258;
    wire N__10255;
    wire N__10252;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10198;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10186;
    wire N__10183;
    wire N__10182;
    wire N__10179;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10171;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10156;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10135;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10125;
    wire N__10122;
    wire N__10117;
    wire N__10116;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10104;
    wire N__10099;
    wire N__10096;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10086;
    wire N__10081;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10038;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10026;
    wire N__10025;
    wire N__10024;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__10005;
    wire N__10002;
    wire N__9999;
    wire N__9996;
    wire N__9991;
    wire N__9988;
    wire N__9985;
    wire N__9980;
    wire N__9973;
    wire N__9970;
    wire N__9967;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9943;
    wire N__9942;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9924;
    wire N__9921;
    wire N__9918;
    wire N__9917;
    wire N__9916;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9900;
    wire N__9897;
    wire N__9892;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9874;
    wire N__9871;
    wire N__9868;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9856;
    wire N__9853;
    wire N__9850;
    wire N__9849;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9826;
    wire N__9825;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9798;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9774;
    wire N__9771;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9744;
    wire N__9741;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9714;
    wire N__9711;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9681;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9657;
    wire N__9654;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9627;
    wire N__9624;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9597;
    wire N__9594;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9574;
    wire N__9571;
    wire N__9568;
    wire N__9567;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9537;
    wire N__9534;
    wire N__9531;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9516;
    wire N__9511;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire N__9492;
    wire N__9487;
    wire N__9484;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9472;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9460;
    wire N__9457;
    wire N__9454;
    wire N__9451;
    wire N__9448;
    wire N__9445;
    wire N__9444;
    wire N__9439;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9402;
    wire N__9401;
    wire N__9394;
    wire N__9393;
    wire N__9390;
    wire N__9387;
    wire N__9382;
    wire N__9381;
    wire N__9380;
    wire N__9379;
    wire N__9376;
    wire N__9375;
    wire N__9374;
    wire N__9367;
    wire N__9364;
    wire N__9359;
    wire N__9356;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9327;
    wire N__9326;
    wire N__9319;
    wire N__9316;
    wire N__9315;
    wire N__9312;
    wire N__9311;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9292;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9282;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9270;
    wire N__9267;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9234;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9138;
    wire N__9137;
    wire N__9130;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9108;
    wire N__9107;
    wire N__9106;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9066;
    wire N__9065;
    wire N__9060;
    wire N__9057;
    wire N__9056;
    wire N__9055;
    wire N__9054;
    wire N__9049;
    wire N__9048;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9030;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8968;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8952;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8928;
    wire N__8927;
    wire N__8926;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8863;
    wire N__8860;
    wire N__8859;
    wire N__8856;
    wire N__8855;
    wire N__8854;
    wire N__8845;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8817;
    wire N__8816;
    wire N__8813;
    wire N__8808;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8784;
    wire N__8783;
    wire N__8782;
    wire N__8781;
    wire N__8778;
    wire N__8773;
    wire N__8768;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8749;
    wire N__8748;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8727;
    wire N__8724;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8704;
    wire N__8701;
    wire N__8698;
    wire N__8697;
    wire N__8694;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8674;
    wire N__8671;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8649;
    wire N__8644;
    wire N__8641;
    wire N__8638;
    wire N__8635;
    wire N__8634;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8619;
    wire N__8614;
    wire N__8611;
    wire N__8608;
    wire N__8607;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8592;
    wire N__8587;
    wire N__8584;
    wire N__8581;
    wire N__8580;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8565;
    wire N__8560;
    wire N__8557;
    wire N__8556;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8535;
    wire N__8532;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8517;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8502;
    wire N__8497;
    wire N__8496;
    wire N__8495;
    wire N__8494;
    wire N__8485;
    wire N__8482;
    wire N__8481;
    wire N__8480;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8373;
    wire N__8372;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8280;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8230;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8139;
    wire N__8138;
    wire N__8135;
    wire N__8130;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8098;
    wire N__8095;
    wire N__8092;
    wire N__8089;
    wire N__8088;
    wire N__8083;
    wire N__8080;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8070;
    wire N__8067;
    wire N__8066;
    wire N__8059;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8040;
    wire N__8039;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8027;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8011;
    wire N__8010;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7990;
    wire N__7987;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7974;
    wire N__7973;
    wire N__7970;
    wire N__7965;
    wire N__7960;
    wire N__7959;
    wire N__7958;
    wire N__7957;
    wire N__7954;
    wire N__7947;
    wire N__7942;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7927;
    wire N__7924;
    wire N__7921;
    wire N__7918;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7908;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7884;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7872;
    wire N__7867;
    wire N__7864;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7852;
    wire N__7849;
    wire N__7848;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7831;
    wire N__7828;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire \latticehx1k_pll_inst.clk ;
    wire clk_in_c;
    wire GNDG0;
    wire VCCG0;
    wire bfn_1_3_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire bfn_1_6_0_;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.N_41_i ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire uart_RXD;
    wire bfn_2_5_0_;
    wire \buart.Z_tx.counter_RNIVE1P1_1 ;
    wire \buart.Z_tx.un1_bitcount_cry_0 ;
    wire \buart.Z_tx.counter_RNIVE1P1_0_1 ;
    wire \buart.Z_tx.un1_bitcount_cry_1 ;
    wire \buart.Z_tx.un1_bitcount_axb_3 ;
    wire \buart.Z_tx.un1_bitcount_cry_2 ;
    wire \buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \ufifo.fifo.fifo_txdata_2 ;
    wire \ufifo.fifo.fifo_txdata_1 ;
    wire \ufifo.sb_ram512x8_inst_RNIKRN11_cascade_ ;
    wire \ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0 ;
    wire utb_txdata_1;
    wire \ufifo.fifo.fifo_txdata_0 ;
    wire \ufifo.fifo.fifo_txdata_6 ;
    wire \ufifo.fifo.fifo_txdata_5 ;
    wire ufifo_utb_txdata_m0_5;
    wire \ufifo.fifo.fifo_txdata_7 ;
    wire ufifo_utb_txdata_m0_7;
    wire ufifo_utb_txdata_m0_6;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire \ufifo.un4_rxDataValidNoEscZ0Z_1_cascade_ ;
    wire \ufifo.rxDataValidNoEscZ0 ;
    wire \ufifo.fifo.fifo_txdata_3 ;
    wire \ufifo.fifo.fifo_txdata_4 ;
    wire \ufifo.utb_txdata_m0_0 ;
    wire utb_txdata_0;
    wire Lab_UT_dk_de_cr_2_reti;
    wire ufifo_utb_txdata_m0_3;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire ufifo_utb_txdata_m0_4;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \Lab_UT.scdp.byteToEncrypt_7 ;
    wire \Lab_UT.scdp.u2.byteToEncrypt_0 ;
    wire bfn_4_1_0_;
    wire \ufifo.fifo.un1_rdaddr_cry_0 ;
    wire \ufifo.fifo.un1_rdaddr_cry_1 ;
    wire \ufifo.fifo.un1_rdaddr_cry_2 ;
    wire \ufifo.fifo.un1_rdaddr_cry_3 ;
    wire \ufifo.fifo.un1_rdaddr_cry_4 ;
    wire \ufifo.fifo.un1_rdaddr_cry_5 ;
    wire \ufifo.fifo.un1_rdaddr_cry_6 ;
    wire \ufifo.fifo.un1_rdaddr_cry_7 ;
    wire bfn_4_2_0_;
    wire bfn_4_3_0_;
    wire \ufifo.fifo.un1_wraddr_cry_0 ;
    wire \ufifo.fifo.un1_wraddr_cry_1 ;
    wire \ufifo.fifo.un1_wraddr_cry_2 ;
    wire \ufifo.fifo.un1_wraddr_cry_3 ;
    wire \ufifo.fifo.un1_wraddr_cry_4 ;
    wire \ufifo.fifo.un1_wraddr_cry_5 ;
    wire \ufifo.fifo.un1_wraddr_cry_6 ;
    wire \ufifo.fifo.un1_wraddr_cry_7 ;
    wire bfn_4_4_0_;
    wire \resetGen.un12_ci_cascade_ ;
    wire \ufifo.fifo.wraddrZ0Z_6 ;
    wire \ufifo.fifo.rdaddrZ0Z_7 ;
    wire \ufifo.fifo.wraddrZ0Z_7 ;
    wire \ufifo.fifo.rdaddrZ0Z_6 ;
    wire \ufifo.fifo.wraddrZ0Z_0 ;
    wire \ufifo.fifo.rdaddrZ0Z_8 ;
    wire \ufifo.fifo.wraddrZ0Z_8 ;
    wire \ufifo.fifo.rdaddrZ0Z_0 ;
    wire \resetGen.reset_countZ0Z_0 ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \Lab_UT.scdp.q_RNI56C1D_0_cascade_ ;
    wire \ufifo.txdataDZ0Z_0 ;
    wire \ufifo.txdataDZ0Z_6 ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire \resetGen.reset_count_2_0_4_cascade_ ;
    wire \resetGen.un12_ci ;
    wire \resetGen.un23_ci ;
    wire \resetGen.escKeyZ0 ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire \Lab_UT.scdp.msBitsi.q_esr_RNIF1M8Z0Z_6 ;
    wire \Lab_UT.scdp.msBitsi.q_esr_RNIQQ8EZ0Z_0 ;
    wire \resetGen.escKey_0Z0Z_0 ;
    wire \Lab_UT.scdp.msBitsi.msBitsD_6 ;
    wire \Lab_UT.scdp.u2.byteToEncryptZ0Z_5 ;
    wire \Lab_UT.scdp.d2eData_5_cascade_ ;
    wire \Lab_UT.scdp.byteToEncrypt_6 ;
    wire \Lab_UT.scdp.N_52_cascade_ ;
    wire \Lab_UT.scdp.msBitsi.msBitsDZ0Z_0 ;
    wire \Lab_UT.scdp.byteToEncrypt_4 ;
    wire \Lab_UT.scdp.b2a0.N_55 ;
    wire \Lab_UT.scdp.d2eData_5 ;
    wire \Lab_UT.scdp.b2a0.N_55_cascade_ ;
    wire \Lab_UT.scdp.a2b.val_0_0Z0Z_3_cascade_ ;
    wire \Lab_UT.scdp.d2eData_3_6 ;
    wire \Lab_UT.scdp.d2eData_3_6_cascade_ ;
    wire \Lab_UT.scdp.u0.byteToDecrypt_6 ;
    wire \ufifo.sb_ram512x8_inst_RNILSN11 ;
    wire \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0_cascade_ ;
    wire ufifo_utb_txdata_sm0_0;
    wire utb_txdata_2;
    wire \ufifo.txdataDZ0Z_1 ;
    wire \Lab_UT.scdp.msBitsi.msBitsD_1 ;
    wire \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8Z0Z_1 ;
    wire \ufifo.txdataDZ0Z_5 ;
    wire \Lab_UT.scdp.u2.sccEldByte_0 ;
    wire \Lab_UT.scdp.msBitsi.msBitsD_2 ;
    wire \Lab_UT.scdp.msBitsi.L4_tx_data_ns_1_2_cascade_ ;
    wire \ufifo.txdataDZ0Z_2 ;
    wire \Lab_UT.scdp.d2eData_3_1_cascade_ ;
    wire \Lab_UT.scdp.q_RNIABC1D_1 ;
    wire \Lab_UT.scdp.u2.byteToEncrypt_1 ;
    wire \Lab_UT.scdp.d2eData_1_cascade_ ;
    wire \Lab_UT.scdp.lsBits_6_cascade_ ;
    wire \Lab_UT.scdp.lsBitsD_1 ;
    wire \Lab_UT.scdp.lsBitsi.lsBitsD_3 ;
    wire \Lab_UT.scdp.byteToEncrypt_3 ;
    wire \Lab_UT.scdp.lsBitsD_6 ;
    wire \Lab_UT.scdp.d2eData_3_2_cascade_ ;
    wire \Lab_UT.scdp.u2.byteToEncrypt_2 ;
    wire \Lab_UT.scdp.d2eData_2 ;
    wire \Lab_UT.scdp.d2eData_1 ;
    wire \Lab_UT.scdp.lsBitsD_2 ;
    wire \Lab_UT.scdp.d2eData_3_1 ;
    wire \Lab_UT.scdp.pinst0.un12_pValidZ0Z_0_cascade_ ;
    wire \Lab_UT.scdp.un12_pValid_cascade_ ;
    wire \Lab_UT.scdp.d2eData_3_0 ;
    wire \Lab_UT.scdp.un12_pValid ;
    wire \Lab_UT.scdp.e2dData_6 ;
    wire \Lab_UT.scdp.q_RNIDHFGA_3 ;
    wire \Lab_UT.scdp.d2eData_3_2 ;
    wire \Lab_UT.scdp.e2dData_2 ;
    wire \Lab_UT.scdp.N_59_i ;
    wire \Lab_UT.scdp.pinst0.un12_pValidZ0Z_1 ;
    wire \Lab_UT.scdp.msBitsi.msBitsD_4 ;
    wire \Lab_UT.scdp.d2eData_3_4 ;
    wire \Lab_UT.scdp.d2eData_3_4_cascade_ ;
    wire \Lab_UT.scdp.q_RNIIAV0D_0_cascade_ ;
    wire \Lab_UT.scdp.msBitsi.q_esr_RNI239EZ0Z_4 ;
    wire \ufifo.txdataDZ0Z_4 ;
    wire \Lab_UT.scdp.d2eData_3_3 ;
    wire \Lab_UT.scdp.pValid_0 ;
    wire \Lab_UT.scdp.d2eData_3_3_cascade_ ;
    wire \Lab_UT.scdp.lsBitsi.q_esr_RNI0TMAZ0Z_3 ;
    wire \Lab_UT.scdp.q_RNIRM8BD_3_cascade_ ;
    wire \ufifo.txdataDZ0Z_3 ;
    wire \Lab_UT.scdp.byteToDecrypt_0 ;
    wire \Lab_UT.scdp.byteToDecrypt_3 ;
    wire \ufifo.fifo.wraddrZ0Z_4 ;
    wire \ufifo.fifo.rdaddrZ0Z_4 ;
    wire \ufifo.fifo.wraddrZ0Z_5 ;
    wire \ufifo.fifo.rdaddrZ0Z_5 ;
    wire \ufifo.fifo.wraddrZ0Z_2 ;
    wire \ufifo.fifo.rdaddrZ0Z_3 ;
    wire \ufifo.fifo.wraddrZ0Z_3 ;
    wire \ufifo.fifo.rdaddrZ0Z_2 ;
    wire \ufifo.fifo.wraddrZ0Z_1 ;
    wire \ufifo.fifo.un1_emptyB_NE_0_cascade_ ;
    wire \ufifo.fifo.rdaddrZ0Z_1 ;
    wire \ufifo.tx_fsm.fifo_txdata_rdy ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \ufifo.fifo.un1_emptyB_NE_2 ;
    wire \ufifo.fifo.un1_emptyB_NE_1 ;
    wire \ufifo.fifo.un1_emptyB_NE_3 ;
    wire \ufifo.fifo.un1_emptyB_NE_4 ;
    wire \ufifo.emptyB_0_cascade_ ;
    wire \ufifo.tx_fsm.cstateZ0Z_1 ;
    wire \ufifo.tx_fsm.N_62_0_cascade_ ;
    wire \ufifo.popFifo ;
    wire rst_i_3_i;
    wire \ufifo.emitcrlf_fsm.cstateZ0Z_0 ;
    wire \buart.Z_rx.bitcountlde_i_o2_0_cascade_ ;
    wire \buart.Z_rx.N_58_cascade_ ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire \buart.Z_rx.N_58 ;
    wire \buart.Z_rx.startbit_cascade_ ;
    wire \buart.Z_rx.ser_clk ;
    wire bfn_5_7_0_;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \buart.Z_rx.N_41_i_1 ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.startbit ;
    wire \buart.Z_rx.N_45 ;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.N_43 ;
    wire \Lab_UT.dk.de_bigL_sxZ0 ;
    wire \Lab_UT.de_bigL_3 ;
    wire \Lab_UT.scctrl.g0_17_N_3LZ0Z3 ;
    wire \Lab_UT.de_bigL_3_cascade_ ;
    wire \Lab_UT.scctrl.g0_17_N_2LZ0Z1 ;
    wire \Lab_UT.de_bigL_0 ;
    wire buart__rx_bitcount_3;
    wire buart__rx_bitcount_0;
    wire buart__rx_bitcount_1;
    wire buart__rx_bitcount_4;
    wire \buart.Z_rx.shifter_0_fast_RNI1CIH1Z0Z_2 ;
    wire \buart.Z_rx.bitcount_es_RNIF6D61Z0Z_4_cascade_ ;
    wire Lab_UT_dk_de_bigD_0;
    wire \Lab_UT.dk.de_bigD_sxZ0 ;
    wire Lab_UT_dk_de_bigD_0_cascade_;
    wire \Lab_UT.dk.de_bigD_1Z0Z_0 ;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_14 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25 ;
    wire \Lab_UT.scdp.prng_lfsr_15 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_3 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10 ;
    wire \Lab_UT.scdp.prng_lfsr_23 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28 ;
    wire \Lab_UT.scdp.prng_lfsr_7 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29 ;
    wire \Lab_UT.scdp.d2eData_3_5 ;
    wire \Lab_UT.scdp.d2eData_3_5_cascade_ ;
    wire \Lab_UT.scdp.e2dData_5 ;
    wire \Lab_UT.scdp.u0.byteToDecrypt_5 ;
    wire \Lab_UT.scdp.u0.byteToDecrypt_7 ;
    wire \Lab_UT.scdp.val_0_3 ;
    wire \Lab_UT.scdp.key1_7 ;
    wire \Lab_UT.scdp.key1_3 ;
    wire \ufifo.txDataValidDZ0 ;
    wire \ufifo.emitcrlf_fsm.cstate_srsts_sn_1 ;
    wire \ufifo.N_57_0_1_cascade_ ;
    wire \ufifo.tx_fsm.cstateZ0Z_4 ;
    wire \ufifo.tx_fsm.N_59_0 ;
    wire buart__tx_uart_busy_0;
    wire \ufifo.emitcrlf_fsm.cstateZ0Z_1 ;
    wire \ufifo.emitcrlf_fsm.cstate_srsts_rn_0_1 ;
    wire \ufifo.tx_fsm.cstateZ0Z_5 ;
    wire \ufifo.crlfdone ;
    wire \ufifo.tx_fsm.N_72_cascade_ ;
    wire \ufifo.cstate_0 ;
    wire \Lab_UT.dk.de_bigEZ0Z_2 ;
    wire \Lab_UT.scctrl.m24_e_4 ;
    wire \Lab_UT.dk.escKey_4_reti_cascade_ ;
    wire \Lab_UT.scctrl.g0_i_a7_1 ;
    wire \Lab_UT.scctrl.g0_i_a3_2_cascade_ ;
    wire \Lab_UT.g0_i_a9_1_3_cascade_ ;
    wire bu_rx_data_rdy_cascade_;
    wire \Lab_UT.scctrl.delay1 ;
    wire \Lab_UT.scctrl.delay2 ;
    wire N_6;
    wire \Lab_UT.scdp.pinst1.un12_pValidZ0Z_1_cascade_ ;
    wire \Lab_UT.un7_pValid ;
    wire \Lab_UT.un1_pValid ;
    wire \Lab_UT.un7_pValid_cascade_ ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_1_0_i_cascade_ ;
    wire \Lab_UT.scctrl.next_state_0_sqmuxa_4Z0Z_0 ;
    wire \Lab_UT.dk.de_bigEZ0Z_1 ;
    wire Lab_UT_dk_de_bigD_6_cascade_;
    wire \Lab_UT.de_bigE_cascade_ ;
    wire \Lab_UT.scdp.N_39_cascade_ ;
    wire \Lab_UT.scdp.a2b.N_50_cascade_ ;
    wire \Lab_UT.scdp.a2b.N_51 ;
    wire bu_rx_data_i_2_5;
    wire \Lab_UT.scctrl.m24_e_5 ;
    wire \Lab_UT.scdp.a2b.N_50 ;
    wire bu_rx_data_3;
    wire \Lab_UT.scdp.a2b.N_53_cascade_ ;
    wire \Lab_UT.scdp.N_39 ;
    wire \Lab_UT.scdp.byteToDecrypt_4 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_6 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsr_next_1_0_cascade_ ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_4 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_11 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_12 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13 ;
    wire \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_g ;
    wire \Lab_UT.scdp.key3_0 ;
    wire buart__rx_bitcount_2;
    wire \buart.Z_rx.bitcount_es_RNIGTPI1Z0Z_3 ;
    wire \Lab_UT.scdp.d2eData_0 ;
    wire \Lab_UT.scdp.lsBitsD_0 ;
    wire \Lab_UT.scdp.lsBits_6 ;
    wire \Lab_UT.scdp.lsBitsD_4 ;
    wire \Lab_UT.scdp.N_48_i ;
    wire \Lab_UT.scdp.N_52 ;
    wire \Lab_UT.scdp.msBitsD_3 ;
    wire buart__tx_uart_busy_0_i;
    wire \buart.Z_tx.N_255 ;
    wire ufifo_utb_txdata_rdy_0;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \Lab_UT.scctrl.delay3 ;
    wire \Lab_UT.scctrl.r4.delay4 ;
    wire \Lab_UT.scdp.u1.byteToDecrypt_2 ;
    wire \Lab_UT.scdp.key1_5 ;
    wire \Lab_UT.scdp.key1_1 ;
    wire \Lab_UT.scdp.key2_5 ;
    wire \Lab_UT.scdp.key3_5 ;
    wire \Lab_UT.scdp.key3_1 ;
    wire \Lab_UT.scdp.key1_0 ;
    wire \Lab_UT.scdp.key2_4 ;
    wire \Lab_UT.scdp.key3_4 ;
    wire \Lab_UT.sccEldByte ;
    wire \Lab_UT.state_ret_6_RNIL97G01_0 ;
    wire \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_iZ0 ;
    wire \Lab_UT.scctrl.un1_state_inv_cascade_ ;
    wire \Lab_UT.scctrl.state_ret_12_RNIUQFKZ0_cascade_ ;
    wire \Lab_UT.state_ret_12_RNIMJCP8_0_cascade_ ;
    wire \Lab_UT.scctrl.delayload ;
    wire \Lab_UT.scctrl.next_state_rst_1_0_cascade_ ;
    wire \Lab_UT.scctrl.un1_state_3_1_reti_cascade_ ;
    wire \Lab_UT.de_bigE_0 ;
    wire \Lab_UT.scctrl.g0_7_1_0 ;
    wire \Lab_UT.scctrl.g2_0_2_cascade_ ;
    wire \Lab_UT.scctrl.g0_2_cascade_ ;
    wire \Lab_UT.scctrl.g0_7_cascade_ ;
    wire \Lab_UT.scctrl.g1_0 ;
    wire \Lab_UT.scctrl.g2_2 ;
    wire \Lab_UT.scctrl.g1 ;
    wire \Lab_UT.sccDnibble1En ;
    wire \Lab_UT.sccDnibble1En_cascade_ ;
    wire \Lab_UT.scdp.u0.sccDnibble1En_0 ;
    wire \Lab_UT.scctrl.next_state_1_sqmuxa_3_0_cascade_ ;
    wire \Lab_UT.scctrl.state_retZ0Z_10 ;
    wire \Lab_UT.scctrl.next_state_1_sqmuxa_3_cascade_ ;
    wire \Lab_UT.scctrl.nibbleInZ0Z1 ;
    wire \Lab_UT.scctrl.N_1_0_i ;
    wire \Lab_UT.scctrl.next_state_1_sqmuxa_3 ;
    wire \Lab_UT.scctrl.un6_sccDecrypt ;
    wire \Lab_UT.de_bigE ;
    wire \Lab_UT.scctrl.next_state_1_i_a5_1_0 ;
    wire \Lab_UT.scctrl.EmsLoaded ;
    wire \Lab_UT.scctrl.EmsLoaded_cascade_ ;
    wire \Lab_UT.sccElsBitsLd_cascade_ ;
    wire \Lab_UT.scdp.sccElsBitsLd_0 ;
    wire \Lab_UT.sccElsBitsLd ;
    wire \Lab_UT.scdp.lsBitsi.lsBitsD_5 ;
    wire Lab_UT_dk_de_cr_12_1_cascade_;
    wire L4_PrintBuf_cascade_;
    wire \Lab_UT.scctrl.N_9_0 ;
    wire bu_rx_data_fast_0;
    wire buart__rx_shifter_0_fast_3;
    wire \Lab_UT.dk.un7_de_hex_xZ0Z0_cascade_ ;
    wire \Lab_UT.dk.un7_de_hex_0_cascade_ ;
    wire \Lab_UT.dk.un7_de_hex_0 ;
    wire \Lab_UT.un4_de_hex_cascade_ ;
    wire buart__rx_shifter_0_fast_1;
    wire buart__rx_shifter_ret_1_fast;
    wire \Lab_UT.scctrl.g0_i_o9_0Z0Z_2 ;
    wire \Lab_UT.dk.un4_de_hexZ0Z_1 ;
    wire bu_rx_data_i_3_4;
    wire bu_rx_data_5;
    wire bu_rx_data_4;
    wire bu_rx_data_i_2_6;
    wire \Lab_UT.un1_de_hex_2 ;
    wire \Lab_UT.un1_de_hex_2_cascade_ ;
    wire \Lab_UT.scctrl.g0_i_a9_3_4_cascade_ ;
    wire \Lab_UT.scctrl.g0_i_a9_3_5 ;
    wire \Lab_UT.scctrl.next_state_1_0_a5_2_out_cascade_ ;
    wire \Lab_UT.scctrl.N_222_1 ;
    wire \Lab_UT.scctrl.next_state_3_sqmuxa_0 ;
    wire \Lab_UT.scdp.a2b.g1_1_a3_0Z0Z_0 ;
    wire \Lab_UT.scdp.key0_0 ;
    wire \Lab_UT.scdp.key0_2 ;
    wire \Lab_UT.scdp.key1_4 ;
    wire \Lab_UT.state_ret_13_RNIQ72741_0 ;
    wire \Lab_UT.scdp.key1_6 ;
    wire \Lab_UT.scctrl.next_state77_cascade_ ;
    wire \Lab_UT.scctrl.next_state_3_sqmuxa ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_0_cascade_ ;
    wire \Lab_UT.scctrl.next_state77 ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_cascade_ ;
    wire \Lab_UT.scctrl.next_state77_2 ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz_4 ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz ;
    wire \Lab_UT.scctrl.next_state76 ;
    wire \Lab_UT.scdp.key2_3 ;
    wire \Lab_UT.scdp.key2_6 ;
    wire \Lab_UT.state_ret_14_RNI416G41_0 ;
    wire \Lab_UT.scdp.key3_6 ;
    wire \Lab_UT.scdp.key3_2 ;
    wire \Lab_UT.state_2_RNI44QH41_0_2 ;
    wire \Lab_UT.scdp.key2_7 ;
    wire \Lab_UT.state_2_RNIF0RJ41_0_2 ;
    wire \Lab_UT.scdp.key3_3 ;
    wire \Lab_UT.state_ret_13_RNIHUNI41_0 ;
    wire \Lab_UT.state_ret_13_RNIHUNI41_0_cascade_ ;
    wire \Lab_UT.scdp.key1_2 ;
    wire \Lab_UT.sccDecrypt_0 ;
    wire \Lab_UT.state_ret_12_RNIMJCP8_0 ;
    wire \Lab_UT.sccDnibble2En_cascade_ ;
    wire resetGen_rst_0_iso;
    wire \Lab_UT.scdp.u1.sccDnibble2En_0 ;
    wire \Lab_UT.scdp.N_37 ;
    wire \Lab_UT.sccDnibble2En ;
    wire \Lab_UT.scdp.byteToDecrypt_1 ;
    wire CONSTANT_ONE_NET;
    wire \Lab_UT.scctrl.g0_i_a9_0_1_cascade_ ;
    wire \Lab_UT.scctrl.g0_i_a9_1 ;
    wire \Lab_UT.scctrl.N_12_cascade_ ;
    wire \Lab_UT.scctrl.g0_i_2 ;
    wire \Lab_UT.scctrl.G_23_0_a9_0_0 ;
    wire \Lab_UT.scctrl.g0_i_a10_2_1_cascade_ ;
    wire \Lab_UT.scctrl.G_23_0_2 ;
    wire \Lab_UT.scctrl.N_2ctr ;
    wire \Lab_UT.scctrl.g0_i_0 ;
    wire \Lab_UT.scctrl.g0_i_4 ;
    wire \Lab_UT.scctrl.N_10 ;
    wire \Lab_UT.scctrl.G_23_0_a9_4_2_cascade_ ;
    wire \Lab_UT.scctrl.G_23_0_3 ;
    wire \Lab_UT.scctrl.G_23_0_a9_3_1 ;
    wire \Lab_UT.scctrl.G_23_0_4 ;
    wire \Lab_UT.scctrl.G_23_0_3_cascade_ ;
    wire \Lab_UT.scctrl.N_3ctr ;
    wire \Lab_UT.scctrl.g0_i_a7_2_0 ;
    wire \Lab_UT.scctrl.next_state_1_i_a5_4_0_0 ;
    wire \Lab_UT.scctrl.N_8_0 ;
    wire \Lab_UT.scctrl.g0_0_i_2_cascade_ ;
    wire \Lab_UT.scctrl.state_i_3_fast_0 ;
    wire \Lab_UT.scctrl.g0_i_1_1_0 ;
    wire \Lab_UT.scdp.a2b.N_6_0 ;
    wire \Lab_UT.scctrl.g0_14_mb_rn_0 ;
    wire \Lab_UT.scctrl.g0_0_i_1_cascade_ ;
    wire \Lab_UT.scctrl.N_7_2 ;
    wire \Lab_UT.scctrl.state_i_3_fast_2 ;
    wire \Lab_UT.scctrl.next_state_1_0_a5_0_0_3 ;
    wire N_127_i_i_1_cascade_;
    wire \Lab_UT.scctrl.N_11_0 ;
    wire \Lab_UT.N_166_0_0 ;
    wire \Lab_UT.scctrl.N_127_i_i_3 ;
    wire \Lab_UT.g1_i_a4_0_2_cascade_ ;
    wire \Lab_UT.next_state_3 ;
    wire \Lab_UT.g0_3_a3_0_4_cascade_ ;
    wire \Lab_UT.scctrl.g0_8_0 ;
    wire \Lab_UT.scdp.a2b.g1_1_o2_0Z0Z_0 ;
    wire \Lab_UT.scdp.a2b.N_6_1_cascade_ ;
    wire \Lab_UT.scdp.a2b.g0_3_a3_0Z0Z_3 ;
    wire \Lab_UT.N_190 ;
    wire \Lab_UT.scctrl.N_6_3_0 ;
    wire \Lab_UT.scctrl.g0_1_1_cascade_ ;
    wire \Lab_UT.scctrl.g0_2_0 ;
    wire \Lab_UT.scctrl.N_12_0 ;
    wire \Lab_UT.scctrl.g0_i_1_0 ;
    wire \Lab_UT.scctrl.g0_i_3_0_cascade_ ;
    wire \Lab_UT.scctrl.un6_sccDecrypt_0 ;
    wire \Lab_UT.scctrl.g1_1_0_cascade_ ;
    wire \Lab_UT.scctrl.g2_0 ;
    wire \Lab_UT.scctrl.g0_1_2_cascade_ ;
    wire \Lab_UT.scctrl.next_state_rst_1_3_1_cascade_ ;
    wire \Lab_UT.next_state_rst_1_3 ;
    wire \Lab_UT.next_state_rst_1_3_cascade_ ;
    wire \Lab_UT.scctrl.N_166_0 ;
    wire \Lab_UT.scctrl.next_state_rst_1_cascade_ ;
    wire led_c_2;
    wire \Lab_UT.scctrl.g0_17_N_4LZ0Z5 ;
    wire \Lab_UT.scctrl.next_state_rst_0_3_N_6_1_cascade_ ;
    wire \Lab_UT.scctrl.g0_i_2_0_cascade_ ;
    wire \Lab_UT.scctrl.next_state_rst_0 ;
    wire \Lab_UT.scctrl.g0_i_2_0 ;
    wire \Lab_UT.scctrl.next_state_rst_0_3_N_6_1 ;
    wire \Lab_UT.g0_3_0 ;
    wire \Lab_UT.scctrl.g0_i_a8_3_0 ;
    wire \Lab_UT.scctrl.N_6_3 ;
    wire \Lab_UT.scctrl.g0_i_1_1_cascade_ ;
    wire \Lab_UT.scctrl.next_state_1_0_1_3_cascade_ ;
    wire \Lab_UT.scctrl.next_state75 ;
    wire \Lab_UT.scctrl.N_7_1 ;
    wire \Lab_UT.scctrl.N_223_2 ;
    wire \Lab_UT.scctrl.next_state73 ;
    wire \Lab_UT.scctrl.next_state73_cascade_ ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i ;
    wire \Lab_UT.state_ret_3_RNII68F41_0_cascade_ ;
    wire \Lab_UT.scdp.key2_0 ;
    wire \Lab_UT.scdp.key2_1 ;
    wire \Lab_UT.state_ret_3_RNII68F41_0 ;
    wire \Lab_UT.scdp.key2_2 ;
    wire bu_rx_data_i_3_1;
    wire \Lab_UT.scdp.key0_5 ;
    wire \Lab_UT.scdp.a2b.N_53 ;
    wire bu_rx_data_1;
    wire bu_rx_data_2;
    wire \Lab_UT.scdp.binValD_2 ;
    wire \Lab_UT.scdp.key0_6 ;
    wire \Lab_UT.scdp.binValD_0 ;
    wire \Lab_UT.scdp.key0_4 ;
    wire \Lab_UT.state_ret_RNIUV0941_0 ;
    wire \Lab_UT.scdp.key0_7 ;
    wire \Lab_UT.scdp.binValD_1 ;
    wire \Lab_UT.scdp.key0_1 ;
    wire \Lab_UT.scdp.binValD_3 ;
    wire \Lab_UT.scdp.binVal_ValidD ;
    wire \Lab_UT.state_0_RNIKFK051_0_1 ;
    wire \Lab_UT.scdp.key0_3 ;
    wire \Lab_UT.scctrl.next_state74 ;
    wire G_23_0_0;
    wire \Lab_UT.scctrl.N_12_1 ;
    wire \Lab_UT.scctrl.N_5_0 ;
    wire \Lab_UT.scctrl.g0_0_i_a8_3_1_0 ;
    wire \Lab_UT.scctrl.g0_0_i_a8_2_1_0_cascade_ ;
    wire \Lab_UT.scctrl.g0_0_i_3_0_cascade_ ;
    wire \Lab_UT.scctrl.N_13 ;
    wire \Lab_UT.scctrl.g0_i_1 ;
    wire \Lab_UT.scctrl.g0_0_i_2 ;
    wire \Lab_UT.scctrl.g0_16_mb_sn ;
    wire \Lab_UT.scctrl.g0_16_mb_rn_0 ;
    wire \Lab_UT.scctrl.g0_0_i_3_0 ;
    wire Lab_UT_dk_de_cr_12_1;
    wire \ufifo.emptyB_0 ;
    wire bu_rx_data_0;
    wire \ufifo.tx_fsm.N_60_0 ;
    wire \Lab_UT.scctrl.N_127_i_i_a6_0_0 ;
    wire \Lab_UT.scctrl.N_11 ;
    wire \Lab_UT.scctrl.G_21_i_a7_1_1 ;
    wire \Lab_UT.m61_i_a2_2 ;
    wire \Lab_UT.scctrl.g0_0_i_0_0 ;
    wire \Lab_UT.N_5_cascade_ ;
    wire \Lab_UT.g0_i_5 ;
    wire \Lab_UT.scctrl.g0_14_mb_sn ;
    wire \Lab_UT.scctrl.g0_0_i_1_1 ;
    wire \Lab_UT.scctrl.N_14 ;
    wire \Lab_UT.scdp.a2b.g0_iZ0Z_4 ;
    wire \Lab_UT.N_5 ;
    wire \Lab_UT.scdp.a2b.g0_iZ0Z_8_cascade_ ;
    wire \Lab_UT.scdp.a2b.g0_3_a3_6 ;
    wire \Lab_UT.de_cr_2 ;
    wire \Lab_UT.de_cr_6_0 ;
    wire \Lab_UT.g0_i_a5_1_3_cascade_ ;
    wire \Lab_UT.scdp.a2b.N_9_1 ;
    wire \Lab_UT.scdp.a2b.g1_1_0_1 ;
    wire \Lab_UT.scctrl.g0_1_3_1 ;
    wire \Lab_UT.scctrl.N_127_i_i_o6_0_1_cascade_ ;
    wire \Lab_UT.scctrl.N_127_i_i_a6_1 ;
    wire \Lab_UT.scctrl.N_190_0_0 ;
    wire \Lab_UT.next_state_rst_0_5 ;
    wire \Lab_UT.scdp.a2b.N_6_4 ;
    wire \Lab_UT.state_ret_8_rep1_RNIHA8U3 ;
    wire \Lab_UT.N_182 ;
    wire \Lab_UT.scdp.a2b.g0_iZ0Z_9 ;
    wire \Lab_UT.state_2_RNI3PVB9_2 ;
    wire \Lab_UT.scctrl.N_182_0 ;
    wire \Lab_UT.scctrl.N_166_0_1 ;
    wire bu_rx_data_0_rep1;
    wire \Lab_UT.scctrl.next_state_1_i_o2_0_d_1_cascade_ ;
    wire buart__rx_shifter_0_fast_2;
    wire \Lab_UT.scctrl.next_state_rst_0_3_N_5L8Z0Z_1_cascade_ ;
    wire Lab_UT_dk_de_bigD_6;
    wire shifter_0_fast_RNI639J4_2;
    wire \Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433_cascade_ ;
    wire \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0 ;
    wire \Lab_UT.de_bigD ;
    wire \Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433 ;
    wire \Lab_UT.de_bigL ;
    wire \Lab_UT.scctrl.next_state_1_i_o2_0_d_1 ;
    wire \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0Z_2 ;
    wire bu_rx_data_6;
    wire bu_rx_data_7;
    wire resetGen_escKey_4;
    wire N_41_i_g;
    wire \Lab_UT.scctrl.g0_2_1 ;
    wire \Lab_UT.scctrl.next_state_rst_0_3_N_6_0 ;
    wire \Lab_UT.scctrl.g1_0_0_cascade_ ;
    wire \Lab_UT.scctrl.g0_1_3 ;
    wire \Lab_UT.scctrl.g0_1_0_0 ;
    wire rst_i_3_rep2;
    wire \Lab_UT.state_ret_8_rep1_RNIJDTUE_1 ;
    wire \Lab_UT.scctrl.next_state_rst_0_5_0_cascade_ ;
    wire \Lab_UT.scctrl.stateZ0Z_3 ;
    wire rst_i_3_rep1;
    wire \Lab_UT.scctrl.g0_i_a8_1 ;
    wire \Lab_UT.scctrl.g0_i_0_0 ;
    wire \Lab_UT.scctrl.g0_7_3 ;
    wire \Lab_UT.scctrl.g0_7_2 ;
    wire \Lab_UT.scctrl.g2_cascade_ ;
    wire \Lab_UT.scctrl.g1_1 ;
    wire \Lab_UT.scctrl.g0_1_0 ;
    wire \Lab_UT.scctrl.N_222i_cascade_ ;
    wire \Lab_UT.scctrl.N_223_1_reti ;
    wire \Lab_UT.scctrl.next_state_rst_2 ;
    wire \Lab_UT.scctrl.N_223_2_reti ;
    wire \Lab_UT.next_state_rst_2_0 ;
    wire \Lab_UT.scctrl.g0_i_3 ;
    wire \Lab_UT.scctrl.N_8 ;
    wire \Lab_UT.scctrl.g0_i_4_0_cascade_ ;
    wire led_c_0;
    wire \Lab_UT.scctrl.N_8_1 ;
    wire \Lab_UT.scctrl.N_8_3 ;
    wire \Lab_UT.scctrl.g0_18_1_cascade_ ;
    wire \Lab_UT.scctrl.next_stateZ0Z_2 ;
    wire \Lab_UT.scctrl.next_stateZ0Z_2_cascade_ ;
    wire \Lab_UT.scctrl.N_6_2 ;
    wire \Lab_UT.scctrl.g0_i_3_1 ;
    wire next_state_1;
    wire \Lab_UT.scctrl.g0_i_m4_1_1 ;
    wire \Lab_UT.scctrl.N_9 ;
    wire \Lab_UT.scctrl.g1_i_a7_1 ;
    wire \Lab_UT.scctrl.next_state_0_3 ;
    wire \Lab_UT.scctrl.next_state_1_0_3 ;
    wire \Lab_UT.scctrl.next_state_i_3_cascade_ ;
    wire \Lab_UT.scctrl.next_state71 ;
    wire \Lab_UT.scctrl.next_state72 ;
    wire \Lab_UT.scctrl.g4_1 ;
    wire \Lab_UT.sccEmsBitsSl ;
    wire \Lab_UT.scctrl.g2 ;
    wire \Lab_UT.scctrl.next_state_rst_3 ;
    wire resetGen_rst_0_iso_g;
    wire \Lab_UT.scctrl.g0_0_i_a8_0_1_cascade_ ;
    wire \Lab_UT.scctrl.N_20 ;
    wire \Lab_UT.scctrl.G_38_0_a3_0_4_cascade_ ;
    wire \Lab_UT.scctrl.next_stateZ0Z_0 ;
    wire \Lab_UT.scctrl.G_38_0_1_cascade_ ;
    wire \Lab_UT.scctrl.N_7_0 ;
    wire \Lab_UT.scctrl.g0_0_i_0 ;
    wire \Lab_UT.scdp.a2b.g0_i_a9_1 ;
    wire \Lab_UT.scdp.a2b.g0_iZ0Z_1_cascade_ ;
    wire \Lab_UT.scdp.a2b.g0_iZ0Z_2 ;
    wire \Lab_UT.scctrl.g0_7_a13_1_1_cascade_ ;
    wire \Lab_UT.scctrl.N_7_cascade_ ;
    wire \Lab_UT.scctrl.g0_6 ;
    wire rst;
    wire \Lab_UT.scctrl.g1_i_a7_2Z0Z_3 ;
    wire \Lab_UT.scctrl.N_10_1_cascade_ ;
    wire \Lab_UT.scctrl.g1_i_2 ;
    wire \Lab_UT.scctrl.N_7_4 ;
    wire \Lab_UT.un1_de_hex ;
    wire \Lab_UT.scctrl.G_21_i_a7_0 ;
    wire \Lab_UT.un4_de_hex ;
    wire \Lab_UT.scctrl.N_11_1 ;
    wire \Lab_UT.scctrl.N_12_2 ;
    wire \Lab_UT.scctrl.G_24_i_a4_1_cascade_ ;
    wire \Lab_UT.scctrl.G_21_i_a7_0_1 ;
    wire \Lab_UT.scctrl.N_9_2 ;
    wire \Lab_UT.scctrl.G_21_i_2 ;
    wire \Lab_UT.scctrl.N_8_2 ;
    wire \Lab_UT.state_i_3_0_rep1 ;
    wire \Lab_UT.state_i_3_2_rep1 ;
    wire \Lab_UT.scctrl.g0_1_4_1 ;
    wire \Lab_UT.scctrl.g0_i_a7_0_1_cascade_ ;
    wire \Lab_UT.de_hex_0 ;
    wire \Lab_UT.scctrl.N_10_0 ;
    wire \Lab_UT.un1_state_3_1 ;
    wire L4_PrintBuf;
    wire \Lab_UT.scctrl.m26_i_o4_1_2 ;
    wire \Lab_UT.scctrl.G_24_i_o3_0_0_cascade_ ;
    wire bu_rx_data_rdy;
    wire \Lab_UT.scctrl.N_6_5_cascade_ ;
    wire \Lab_UT.scctrl.N_5_2 ;
    wire \Lab_UT.scctrl.N_8_4 ;
    wire \Lab_UT.scctrl.N_4ctr ;
    wire \Lab_UT.scctrl.G_23_0_a9_1 ;
    wire \Lab_UT.state_i_3_1 ;
    wire \Lab_UT.scctrl.g0_i_a8_4_1 ;
    wire \Lab_UT.scctrl.next_state_0_2 ;
    wire rst_i_3;
    wire Lab_UT_scctrl_N_221_0;
    wire \Lab_UT.scctrl.G_21_i_0 ;
    wire \Lab_UT.state_i_3_2 ;
    wire \Lab_UT.state_2 ;
    wire \Lab_UT.state_0 ;
    wire \Lab_UT.scctrl.g0_i_7_1 ;
    wire rst_i_3_reti;
    wire clk_g;
    wire \Lab_UT.scctrl.g2_1 ;
    wire \Lab_UT.state_i_3_2_rep2 ;
    wire \Lab_UT.state_i_3_3 ;
    wire \Lab_UT.scctrl.state_i_3_0_rep2 ;
    wire rst_i_3_fast;
    wire \Lab_UT.scctrl.g1_i_0 ;
    wire \Lab_UT.state_i_3_0 ;
    wire \Lab_UT.scctrl.g0_0_i_a8_3_1 ;
    wire \Lab_UT.state_1 ;
    wire \Lab_UT.scctrl.state_1_RNO_3Z0Z_0 ;
    wire \Lab_UT.scctrl.N_13_0 ;
    wire \Lab_UT.N_191 ;
    wire \Lab_UT.scctrl.G_24_i_a4_0_1 ;
    wire \Lab_UT.next_state_1_0_0_3 ;
    wire \Lab_UT.scctrl.N_10_2 ;
    wire \Lab_UT.N_169_0 ;
    wire \Lab_UT.scctrl.N_223_1 ;
    wire led_c_4;
    wire _gnd_net_;

    defparam \ufifo.fifo.sb_ram512x8_inst_physical .WRITE_MODE=1;
    defparam \ufifo.fifo.sb_ram512x8_inst_physical .READ_MODE=1;
    SB_RAM40_4K \ufifo.fifo.sb_ram512x8_inst_physical  (
            .RDATA({dangling_wire_0,\ufifo.fifo.fifo_txdata_7 ,dangling_wire_1,\ufifo.fifo.fifo_txdata_6 ,dangling_wire_2,\ufifo.fifo.fifo_txdata_5 ,dangling_wire_3,\ufifo.fifo.fifo_txdata_4 ,dangling_wire_4,\ufifo.fifo.fifo_txdata_3 ,dangling_wire_5,\ufifo.fifo.fifo_txdata_2 ,dangling_wire_6,\ufifo.fifo.fifo_txdata_1 ,dangling_wire_7,\ufifo.fifo.fifo_txdata_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__8587,N__8704,N__8644,N__9721,N__9781,N__9664,N__9604,N__9544,N__8527}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__8560,N__8674,N__8734,N__9751,N__9808,N__9634,N__9691,N__9574,N__8614}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__8827,dangling_wire_31,N__8983,dangling_wire_32,N__9415,dangling_wire_33,N__9868,dangling_wire_34,N__9193,dangling_wire_35,N__9010,dangling_wire_36,N__8833}),
            .RCLKE(N__10025),
            .RCLK(N__22671),
            .RE(N__10026),
            .WCLKE(N__11091),
            .WCLK(N__22670),
            .WE(N__11092));
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\latticehx1k_pll_inst.clk ),
            .REFERENCECLK(N__7825),
            .RESETB(N__13966),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    IO_PAD led_obuf_4_iopad (
            .OE(N__23195),
            .DIN(N__23194),
            .DOUT(N__23193),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__23195),
            .PADOUT(N__23194),
            .PADIN(N__23193),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21214),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_1_iopad (
            .OE(N__23186),
            .DIN(N__23185),
            .DOUT(N__23184),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__23186),
            .PADOUT(N__23185),
            .PADIN(N__23184),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17807),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_3_iopad (
            .OE(N__23177),
            .DIN(N__23176),
            .DOUT(N__23175),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__23177),
            .PADOUT(N__23176),
            .PADIN(N__23175),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_0_iopad (
            .OE(N__23168),
            .DIN(N__23167),
            .DOUT(N__23166),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__23168),
            .PADOUT(N__23167),
            .PADIN(N__23166),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17808),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__23159),
            .DIN(N__23158),
            .DOUT(N__23157),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__23159),
            .PADOUT(N__23158),
            .PADIN(N__23157),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__22662),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__23150),
            .DIN(N__23149),
            .DOUT(N__23148),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__23150),
            .PADOUT(N__23149),
            .PADIN(N__23148),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__23141),
            .DIN(N__23140),
            .DOUT(N__23139),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__23141),
            .PADOUT(N__23140),
            .PADIN(N__23139),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__23132),
            .DIN(N__23131),
            .DOUT(N__23130),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__23132),
            .PADOUT(N__23131),
            .PADIN(N__23130),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8107),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__23123),
            .DIN(N__23122),
            .DOUT(N__23121),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__23123),
            .PADOUT(N__23122),
            .PADIN(N__23121),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_2_iopad (
            .OE(N__23114),
            .DIN(N__23113),
            .DOUT(N__23112),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__23114),
            .PADOUT(N__23113),
            .PADIN(N__23112),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14672),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__5743 (
            .O(N__23095),
            .I(N__23083));
    CascadeMux I__5742 (
            .O(N__23094),
            .I(N__23080));
    InMux I__5741 (
            .O(N__23093),
            .I(N__23069));
    InMux I__5740 (
            .O(N__23092),
            .I(N__23066));
    InMux I__5739 (
            .O(N__23091),
            .I(N__23057));
    InMux I__5738 (
            .O(N__23090),
            .I(N__23057));
    CascadeMux I__5737 (
            .O(N__23089),
            .I(N__23054));
    InMux I__5736 (
            .O(N__23088),
            .I(N__23048));
    InMux I__5735 (
            .O(N__23087),
            .I(N__23045));
    InMux I__5734 (
            .O(N__23086),
            .I(N__23042));
    InMux I__5733 (
            .O(N__23083),
            .I(N__23039));
    InMux I__5732 (
            .O(N__23080),
            .I(N__23036));
    InMux I__5731 (
            .O(N__23079),
            .I(N__23031));
    InMux I__5730 (
            .O(N__23078),
            .I(N__23031));
    InMux I__5729 (
            .O(N__23077),
            .I(N__23026));
    InMux I__5728 (
            .O(N__23076),
            .I(N__23026));
    CascadeMux I__5727 (
            .O(N__23075),
            .I(N__23023));
    InMux I__5726 (
            .O(N__23074),
            .I(N__23015));
    CascadeMux I__5725 (
            .O(N__23073),
            .I(N__23012));
    CascadeMux I__5724 (
            .O(N__23072),
            .I(N__23008));
    LocalMux I__5723 (
            .O(N__23069),
            .I(N__23003));
    LocalMux I__5722 (
            .O(N__23066),
            .I(N__23003));
    InMux I__5721 (
            .O(N__23065),
            .I(N__22998));
    CascadeMux I__5720 (
            .O(N__23064),
            .I(N__22995));
    InMux I__5719 (
            .O(N__23063),
            .I(N__22988));
    InMux I__5718 (
            .O(N__23062),
            .I(N__22988));
    LocalMux I__5717 (
            .O(N__23057),
            .I(N__22985));
    InMux I__5716 (
            .O(N__23054),
            .I(N__22976));
    InMux I__5715 (
            .O(N__23053),
            .I(N__22976));
    InMux I__5714 (
            .O(N__23052),
            .I(N__22976));
    InMux I__5713 (
            .O(N__23051),
            .I(N__22976));
    LocalMux I__5712 (
            .O(N__23048),
            .I(N__22971));
    LocalMux I__5711 (
            .O(N__23045),
            .I(N__22971));
    LocalMux I__5710 (
            .O(N__23042),
            .I(N__22968));
    LocalMux I__5709 (
            .O(N__23039),
            .I(N__22961));
    LocalMux I__5708 (
            .O(N__23036),
            .I(N__22961));
    LocalMux I__5707 (
            .O(N__23031),
            .I(N__22961));
    LocalMux I__5706 (
            .O(N__23026),
            .I(N__22958));
    InMux I__5705 (
            .O(N__23023),
            .I(N__22950));
    InMux I__5704 (
            .O(N__23022),
            .I(N__22950));
    InMux I__5703 (
            .O(N__23021),
            .I(N__22947));
    InMux I__5702 (
            .O(N__23020),
            .I(N__22944));
    CascadeMux I__5701 (
            .O(N__23019),
            .I(N__22941));
    InMux I__5700 (
            .O(N__23018),
            .I(N__22938));
    LocalMux I__5699 (
            .O(N__23015),
            .I(N__22935));
    InMux I__5698 (
            .O(N__23012),
            .I(N__22932));
    InMux I__5697 (
            .O(N__23011),
            .I(N__22927));
    InMux I__5696 (
            .O(N__23008),
            .I(N__22927));
    IoSpan4Mux I__5695 (
            .O(N__23003),
            .I(N__22924));
    InMux I__5694 (
            .O(N__23002),
            .I(N__22921));
    InMux I__5693 (
            .O(N__23001),
            .I(N__22916));
    LocalMux I__5692 (
            .O(N__22998),
            .I(N__22913));
    InMux I__5691 (
            .O(N__22995),
            .I(N__22910));
    InMux I__5690 (
            .O(N__22994),
            .I(N__22907));
    InMux I__5689 (
            .O(N__22993),
            .I(N__22904));
    LocalMux I__5688 (
            .O(N__22988),
            .I(N__22891));
    Span4Mux_h I__5687 (
            .O(N__22985),
            .I(N__22891));
    LocalMux I__5686 (
            .O(N__22976),
            .I(N__22891));
    Span4Mux_v I__5685 (
            .O(N__22971),
            .I(N__22891));
    Span4Mux_v I__5684 (
            .O(N__22968),
            .I(N__22891));
    Span4Mux_v I__5683 (
            .O(N__22961),
            .I(N__22891));
    Span4Mux_h I__5682 (
            .O(N__22958),
            .I(N__22888));
    InMux I__5681 (
            .O(N__22957),
            .I(N__22881));
    InMux I__5680 (
            .O(N__22956),
            .I(N__22881));
    InMux I__5679 (
            .O(N__22955),
            .I(N__22881));
    LocalMux I__5678 (
            .O(N__22950),
            .I(N__22874));
    LocalMux I__5677 (
            .O(N__22947),
            .I(N__22874));
    LocalMux I__5676 (
            .O(N__22944),
            .I(N__22874));
    InMux I__5675 (
            .O(N__22941),
            .I(N__22871));
    LocalMux I__5674 (
            .O(N__22938),
            .I(N__22866));
    Span4Mux_h I__5673 (
            .O(N__22935),
            .I(N__22866));
    LocalMux I__5672 (
            .O(N__22932),
            .I(N__22863));
    LocalMux I__5671 (
            .O(N__22927),
            .I(N__22860));
    IoSpan4Mux I__5670 (
            .O(N__22924),
            .I(N__22857));
    LocalMux I__5669 (
            .O(N__22921),
            .I(N__22854));
    InMux I__5668 (
            .O(N__22920),
            .I(N__22849));
    InMux I__5667 (
            .O(N__22919),
            .I(N__22849));
    LocalMux I__5666 (
            .O(N__22916),
            .I(N__22846));
    Span4Mux_v I__5665 (
            .O(N__22913),
            .I(N__22835));
    LocalMux I__5664 (
            .O(N__22910),
            .I(N__22835));
    LocalMux I__5663 (
            .O(N__22907),
            .I(N__22835));
    LocalMux I__5662 (
            .O(N__22904),
            .I(N__22835));
    Span4Mux_v I__5661 (
            .O(N__22891),
            .I(N__22835));
    Span4Mux_v I__5660 (
            .O(N__22888),
            .I(N__22828));
    LocalMux I__5659 (
            .O(N__22881),
            .I(N__22828));
    Span4Mux_h I__5658 (
            .O(N__22874),
            .I(N__22828));
    LocalMux I__5657 (
            .O(N__22871),
            .I(N__22817));
    Span4Mux_v I__5656 (
            .O(N__22866),
            .I(N__22817));
    Span4Mux_h I__5655 (
            .O(N__22863),
            .I(N__22817));
    Span4Mux_h I__5654 (
            .O(N__22860),
            .I(N__22817));
    Span4Mux_s1_h I__5653 (
            .O(N__22857),
            .I(N__22817));
    Span12Mux_s1_h I__5652 (
            .O(N__22854),
            .I(N__22814));
    LocalMux I__5651 (
            .O(N__22849),
            .I(\Lab_UT.state_0 ));
    Odrv12 I__5650 (
            .O(N__22846),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__5649 (
            .O(N__22835),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__5648 (
            .O(N__22828),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__5647 (
            .O(N__22817),
            .I(\Lab_UT.state_0 ));
    Odrv12 I__5646 (
            .O(N__22814),
            .I(\Lab_UT.state_0 ));
    CascadeMux I__5645 (
            .O(N__22801),
            .I(N__22798));
    InMux I__5644 (
            .O(N__22798),
            .I(N__22795));
    LocalMux I__5643 (
            .O(N__22795),
            .I(N__22792));
    Odrv4 I__5642 (
            .O(N__22792),
            .I(\Lab_UT.scctrl.g0_i_7_1 ));
    InMux I__5641 (
            .O(N__22789),
            .I(N__22785));
    InMux I__5640 (
            .O(N__22788),
            .I(N__22782));
    LocalMux I__5639 (
            .O(N__22785),
            .I(N__22775));
    LocalMux I__5638 (
            .O(N__22782),
            .I(N__22775));
    InMux I__5637 (
            .O(N__22781),
            .I(N__22772));
    InMux I__5636 (
            .O(N__22780),
            .I(N__22769));
    Span4Mux_v I__5635 (
            .O(N__22775),
            .I(N__22758));
    LocalMux I__5634 (
            .O(N__22772),
            .I(N__22753));
    LocalMux I__5633 (
            .O(N__22769),
            .I(N__22753));
    InMux I__5632 (
            .O(N__22768),
            .I(N__22748));
    InMux I__5631 (
            .O(N__22767),
            .I(N__22748));
    CascadeMux I__5630 (
            .O(N__22766),
            .I(N__22745));
    InMux I__5629 (
            .O(N__22765),
            .I(N__22737));
    InMux I__5628 (
            .O(N__22764),
            .I(N__22737));
    InMux I__5627 (
            .O(N__22763),
            .I(N__22737));
    InMux I__5626 (
            .O(N__22762),
            .I(N__22734));
    InMux I__5625 (
            .O(N__22761),
            .I(N__22731));
    Span4Mux_h I__5624 (
            .O(N__22758),
            .I(N__22724));
    Span4Mux_v I__5623 (
            .O(N__22753),
            .I(N__22724));
    LocalMux I__5622 (
            .O(N__22748),
            .I(N__22724));
    InMux I__5621 (
            .O(N__22745),
            .I(N__22719));
    InMux I__5620 (
            .O(N__22744),
            .I(N__22719));
    LocalMux I__5619 (
            .O(N__22737),
            .I(N__22716));
    LocalMux I__5618 (
            .O(N__22734),
            .I(N__22711));
    LocalMux I__5617 (
            .O(N__22731),
            .I(N__22711));
    Span4Mux_h I__5616 (
            .O(N__22724),
            .I(N__22708));
    LocalMux I__5615 (
            .O(N__22719),
            .I(rst_i_3_reti));
    Odrv12 I__5614 (
            .O(N__22716),
            .I(rst_i_3_reti));
    Odrv12 I__5613 (
            .O(N__22711),
            .I(rst_i_3_reti));
    Odrv4 I__5612 (
            .O(N__22708),
            .I(rst_i_3_reti));
    ClkMux I__5611 (
            .O(N__22699),
            .I(N__22441));
    ClkMux I__5610 (
            .O(N__22698),
            .I(N__22441));
    ClkMux I__5609 (
            .O(N__22697),
            .I(N__22441));
    ClkMux I__5608 (
            .O(N__22696),
            .I(N__22441));
    ClkMux I__5607 (
            .O(N__22695),
            .I(N__22441));
    ClkMux I__5606 (
            .O(N__22694),
            .I(N__22441));
    ClkMux I__5605 (
            .O(N__22693),
            .I(N__22441));
    ClkMux I__5604 (
            .O(N__22692),
            .I(N__22441));
    ClkMux I__5603 (
            .O(N__22691),
            .I(N__22441));
    ClkMux I__5602 (
            .O(N__22690),
            .I(N__22441));
    ClkMux I__5601 (
            .O(N__22689),
            .I(N__22441));
    ClkMux I__5600 (
            .O(N__22688),
            .I(N__22441));
    ClkMux I__5599 (
            .O(N__22687),
            .I(N__22441));
    ClkMux I__5598 (
            .O(N__22686),
            .I(N__22441));
    ClkMux I__5597 (
            .O(N__22685),
            .I(N__22441));
    ClkMux I__5596 (
            .O(N__22684),
            .I(N__22441));
    ClkMux I__5595 (
            .O(N__22683),
            .I(N__22441));
    ClkMux I__5594 (
            .O(N__22682),
            .I(N__22441));
    ClkMux I__5593 (
            .O(N__22681),
            .I(N__22441));
    ClkMux I__5592 (
            .O(N__22680),
            .I(N__22441));
    ClkMux I__5591 (
            .O(N__22679),
            .I(N__22441));
    ClkMux I__5590 (
            .O(N__22678),
            .I(N__22441));
    ClkMux I__5589 (
            .O(N__22677),
            .I(N__22441));
    ClkMux I__5588 (
            .O(N__22676),
            .I(N__22441));
    ClkMux I__5587 (
            .O(N__22675),
            .I(N__22441));
    ClkMux I__5586 (
            .O(N__22674),
            .I(N__22441));
    ClkMux I__5585 (
            .O(N__22673),
            .I(N__22441));
    ClkMux I__5584 (
            .O(N__22672),
            .I(N__22441));
    ClkMux I__5583 (
            .O(N__22671),
            .I(N__22441));
    ClkMux I__5582 (
            .O(N__22670),
            .I(N__22441));
    ClkMux I__5581 (
            .O(N__22669),
            .I(N__22441));
    ClkMux I__5580 (
            .O(N__22668),
            .I(N__22441));
    ClkMux I__5579 (
            .O(N__22667),
            .I(N__22441));
    ClkMux I__5578 (
            .O(N__22666),
            .I(N__22441));
    ClkMux I__5577 (
            .O(N__22665),
            .I(N__22441));
    ClkMux I__5576 (
            .O(N__22664),
            .I(N__22441));
    ClkMux I__5575 (
            .O(N__22663),
            .I(N__22441));
    ClkMux I__5574 (
            .O(N__22662),
            .I(N__22441));
    ClkMux I__5573 (
            .O(N__22661),
            .I(N__22441));
    ClkMux I__5572 (
            .O(N__22660),
            .I(N__22441));
    ClkMux I__5571 (
            .O(N__22659),
            .I(N__22441));
    ClkMux I__5570 (
            .O(N__22658),
            .I(N__22441));
    ClkMux I__5569 (
            .O(N__22657),
            .I(N__22441));
    ClkMux I__5568 (
            .O(N__22656),
            .I(N__22441));
    ClkMux I__5567 (
            .O(N__22655),
            .I(N__22441));
    ClkMux I__5566 (
            .O(N__22654),
            .I(N__22441));
    ClkMux I__5565 (
            .O(N__22653),
            .I(N__22441));
    ClkMux I__5564 (
            .O(N__22652),
            .I(N__22441));
    ClkMux I__5563 (
            .O(N__22651),
            .I(N__22441));
    ClkMux I__5562 (
            .O(N__22650),
            .I(N__22441));
    ClkMux I__5561 (
            .O(N__22649),
            .I(N__22441));
    ClkMux I__5560 (
            .O(N__22648),
            .I(N__22441));
    ClkMux I__5559 (
            .O(N__22647),
            .I(N__22441));
    ClkMux I__5558 (
            .O(N__22646),
            .I(N__22441));
    ClkMux I__5557 (
            .O(N__22645),
            .I(N__22441));
    ClkMux I__5556 (
            .O(N__22644),
            .I(N__22441));
    ClkMux I__5555 (
            .O(N__22643),
            .I(N__22441));
    ClkMux I__5554 (
            .O(N__22642),
            .I(N__22441));
    ClkMux I__5553 (
            .O(N__22641),
            .I(N__22441));
    ClkMux I__5552 (
            .O(N__22640),
            .I(N__22441));
    ClkMux I__5551 (
            .O(N__22639),
            .I(N__22441));
    ClkMux I__5550 (
            .O(N__22638),
            .I(N__22441));
    ClkMux I__5549 (
            .O(N__22637),
            .I(N__22441));
    ClkMux I__5548 (
            .O(N__22636),
            .I(N__22441));
    ClkMux I__5547 (
            .O(N__22635),
            .I(N__22441));
    ClkMux I__5546 (
            .O(N__22634),
            .I(N__22441));
    ClkMux I__5545 (
            .O(N__22633),
            .I(N__22441));
    ClkMux I__5544 (
            .O(N__22632),
            .I(N__22441));
    ClkMux I__5543 (
            .O(N__22631),
            .I(N__22441));
    ClkMux I__5542 (
            .O(N__22630),
            .I(N__22441));
    ClkMux I__5541 (
            .O(N__22629),
            .I(N__22441));
    ClkMux I__5540 (
            .O(N__22628),
            .I(N__22441));
    ClkMux I__5539 (
            .O(N__22627),
            .I(N__22441));
    ClkMux I__5538 (
            .O(N__22626),
            .I(N__22441));
    ClkMux I__5537 (
            .O(N__22625),
            .I(N__22441));
    ClkMux I__5536 (
            .O(N__22624),
            .I(N__22441));
    ClkMux I__5535 (
            .O(N__22623),
            .I(N__22441));
    ClkMux I__5534 (
            .O(N__22622),
            .I(N__22441));
    ClkMux I__5533 (
            .O(N__22621),
            .I(N__22441));
    ClkMux I__5532 (
            .O(N__22620),
            .I(N__22441));
    ClkMux I__5531 (
            .O(N__22619),
            .I(N__22441));
    ClkMux I__5530 (
            .O(N__22618),
            .I(N__22441));
    ClkMux I__5529 (
            .O(N__22617),
            .I(N__22441));
    ClkMux I__5528 (
            .O(N__22616),
            .I(N__22441));
    ClkMux I__5527 (
            .O(N__22615),
            .I(N__22441));
    ClkMux I__5526 (
            .O(N__22614),
            .I(N__22441));
    GlobalMux I__5525 (
            .O(N__22441),
            .I(N__22438));
    gio2CtrlBuf I__5524 (
            .O(N__22438),
            .I(clk_g));
    InMux I__5523 (
            .O(N__22435),
            .I(N__22432));
    LocalMux I__5522 (
            .O(N__22432),
            .I(N__22429));
    Span4Mux_h I__5521 (
            .O(N__22429),
            .I(N__22426));
    Odrv4 I__5520 (
            .O(N__22426),
            .I(\Lab_UT.scctrl.g2_1 ));
    InMux I__5519 (
            .O(N__22423),
            .I(N__22417));
    CascadeMux I__5518 (
            .O(N__22422),
            .I(N__22411));
    InMux I__5517 (
            .O(N__22421),
            .I(N__22408));
    CascadeMux I__5516 (
            .O(N__22420),
            .I(N__22403));
    LocalMux I__5515 (
            .O(N__22417),
            .I(N__22399));
    InMux I__5514 (
            .O(N__22416),
            .I(N__22396));
    InMux I__5513 (
            .O(N__22415),
            .I(N__22393));
    InMux I__5512 (
            .O(N__22414),
            .I(N__22390));
    InMux I__5511 (
            .O(N__22411),
            .I(N__22387));
    LocalMux I__5510 (
            .O(N__22408),
            .I(N__22384));
    InMux I__5509 (
            .O(N__22407),
            .I(N__22379));
    InMux I__5508 (
            .O(N__22406),
            .I(N__22379));
    InMux I__5507 (
            .O(N__22403),
            .I(N__22373));
    InMux I__5506 (
            .O(N__22402),
            .I(N__22373));
    Span12Mux_s3_h I__5505 (
            .O(N__22399),
            .I(N__22370));
    LocalMux I__5504 (
            .O(N__22396),
            .I(N__22365));
    LocalMux I__5503 (
            .O(N__22393),
            .I(N__22365));
    LocalMux I__5502 (
            .O(N__22390),
            .I(N__22360));
    LocalMux I__5501 (
            .O(N__22387),
            .I(N__22360));
    Span4Mux_s3_h I__5500 (
            .O(N__22384),
            .I(N__22355));
    LocalMux I__5499 (
            .O(N__22379),
            .I(N__22355));
    InMux I__5498 (
            .O(N__22378),
            .I(N__22352));
    LocalMux I__5497 (
            .O(N__22373),
            .I(\Lab_UT.state_i_3_2_rep2 ));
    Odrv12 I__5496 (
            .O(N__22370),
            .I(\Lab_UT.state_i_3_2_rep2 ));
    Odrv12 I__5495 (
            .O(N__22365),
            .I(\Lab_UT.state_i_3_2_rep2 ));
    Odrv4 I__5494 (
            .O(N__22360),
            .I(\Lab_UT.state_i_3_2_rep2 ));
    Odrv4 I__5493 (
            .O(N__22355),
            .I(\Lab_UT.state_i_3_2_rep2 ));
    LocalMux I__5492 (
            .O(N__22352),
            .I(\Lab_UT.state_i_3_2_rep2 ));
    CascadeMux I__5491 (
            .O(N__22339),
            .I(N__22336));
    InMux I__5490 (
            .O(N__22336),
            .I(N__22328));
    InMux I__5489 (
            .O(N__22335),
            .I(N__22320));
    InMux I__5488 (
            .O(N__22334),
            .I(N__22316));
    CascadeMux I__5487 (
            .O(N__22333),
            .I(N__22313));
    CascadeMux I__5486 (
            .O(N__22332),
            .I(N__22309));
    CascadeMux I__5485 (
            .O(N__22331),
            .I(N__22306));
    LocalMux I__5484 (
            .O(N__22328),
            .I(N__22298));
    InMux I__5483 (
            .O(N__22327),
            .I(N__22293));
    InMux I__5482 (
            .O(N__22326),
            .I(N__22284));
    InMux I__5481 (
            .O(N__22325),
            .I(N__22284));
    InMux I__5480 (
            .O(N__22324),
            .I(N__22284));
    InMux I__5479 (
            .O(N__22323),
            .I(N__22284));
    LocalMux I__5478 (
            .O(N__22320),
            .I(N__22281));
    InMux I__5477 (
            .O(N__22319),
            .I(N__22278));
    LocalMux I__5476 (
            .O(N__22316),
            .I(N__22275));
    InMux I__5475 (
            .O(N__22313),
            .I(N__22270));
    InMux I__5474 (
            .O(N__22312),
            .I(N__22270));
    InMux I__5473 (
            .O(N__22309),
            .I(N__22263));
    InMux I__5472 (
            .O(N__22306),
            .I(N__22263));
    InMux I__5471 (
            .O(N__22305),
            .I(N__22260));
    CascadeMux I__5470 (
            .O(N__22304),
            .I(N__22254));
    InMux I__5469 (
            .O(N__22303),
            .I(N__22248));
    InMux I__5468 (
            .O(N__22302),
            .I(N__22248));
    InMux I__5467 (
            .O(N__22301),
            .I(N__22245));
    Span4Mux_v I__5466 (
            .O(N__22298),
            .I(N__22242));
    InMux I__5465 (
            .O(N__22297),
            .I(N__22239));
    InMux I__5464 (
            .O(N__22296),
            .I(N__22236));
    LocalMux I__5463 (
            .O(N__22293),
            .I(N__22231));
    LocalMux I__5462 (
            .O(N__22284),
            .I(N__22231));
    Span4Mux_s3_v I__5461 (
            .O(N__22281),
            .I(N__22226));
    LocalMux I__5460 (
            .O(N__22278),
            .I(N__22226));
    Span4Mux_s3_v I__5459 (
            .O(N__22275),
            .I(N__22221));
    LocalMux I__5458 (
            .O(N__22270),
            .I(N__22221));
    InMux I__5457 (
            .O(N__22269),
            .I(N__22216));
    InMux I__5456 (
            .O(N__22268),
            .I(N__22216));
    LocalMux I__5455 (
            .O(N__22263),
            .I(N__22213));
    LocalMux I__5454 (
            .O(N__22260),
            .I(N__22210));
    InMux I__5453 (
            .O(N__22259),
            .I(N__22207));
    InMux I__5452 (
            .O(N__22258),
            .I(N__22202));
    InMux I__5451 (
            .O(N__22257),
            .I(N__22202));
    InMux I__5450 (
            .O(N__22254),
            .I(N__22199));
    InMux I__5449 (
            .O(N__22253),
            .I(N__22196));
    LocalMux I__5448 (
            .O(N__22248),
            .I(N__22193));
    LocalMux I__5447 (
            .O(N__22245),
            .I(N__22187));
    Span4Mux_v I__5446 (
            .O(N__22242),
            .I(N__22184));
    LocalMux I__5445 (
            .O(N__22239),
            .I(N__22177));
    LocalMux I__5444 (
            .O(N__22236),
            .I(N__22177));
    Span4Mux_v I__5443 (
            .O(N__22231),
            .I(N__22177));
    Span4Mux_v I__5442 (
            .O(N__22226),
            .I(N__22172));
    Span4Mux_v I__5441 (
            .O(N__22221),
            .I(N__22172));
    LocalMux I__5440 (
            .O(N__22216),
            .I(N__22169));
    Span4Mux_s2_h I__5439 (
            .O(N__22213),
            .I(N__22160));
    Span4Mux_h I__5438 (
            .O(N__22210),
            .I(N__22160));
    LocalMux I__5437 (
            .O(N__22207),
            .I(N__22160));
    LocalMux I__5436 (
            .O(N__22202),
            .I(N__22160));
    LocalMux I__5435 (
            .O(N__22199),
            .I(N__22153));
    LocalMux I__5434 (
            .O(N__22196),
            .I(N__22153));
    Span4Mux_v I__5433 (
            .O(N__22193),
            .I(N__22153));
    CascadeMux I__5432 (
            .O(N__22192),
            .I(N__22149));
    CascadeMux I__5431 (
            .O(N__22191),
            .I(N__22146));
    CascadeMux I__5430 (
            .O(N__22190),
            .I(N__22143));
    Span4Mux_s2_h I__5429 (
            .O(N__22187),
            .I(N__22140));
    Span4Mux_v I__5428 (
            .O(N__22184),
            .I(N__22135));
    Span4Mux_v I__5427 (
            .O(N__22177),
            .I(N__22135));
    Span4Mux_v I__5426 (
            .O(N__22172),
            .I(N__22130));
    Span4Mux_h I__5425 (
            .O(N__22169),
            .I(N__22130));
    Span4Mux_v I__5424 (
            .O(N__22160),
            .I(N__22125));
    Span4Mux_h I__5423 (
            .O(N__22153),
            .I(N__22125));
    InMux I__5422 (
            .O(N__22152),
            .I(N__22120));
    InMux I__5421 (
            .O(N__22149),
            .I(N__22120));
    InMux I__5420 (
            .O(N__22146),
            .I(N__22115));
    InMux I__5419 (
            .O(N__22143),
            .I(N__22115));
    Odrv4 I__5418 (
            .O(N__22140),
            .I(\Lab_UT.state_i_3_3 ));
    Odrv4 I__5417 (
            .O(N__22135),
            .I(\Lab_UT.state_i_3_3 ));
    Odrv4 I__5416 (
            .O(N__22130),
            .I(\Lab_UT.state_i_3_3 ));
    Odrv4 I__5415 (
            .O(N__22125),
            .I(\Lab_UT.state_i_3_3 ));
    LocalMux I__5414 (
            .O(N__22120),
            .I(\Lab_UT.state_i_3_3 ));
    LocalMux I__5413 (
            .O(N__22115),
            .I(\Lab_UT.state_i_3_3 ));
    CascadeMux I__5412 (
            .O(N__22102),
            .I(N__22097));
    CascadeMux I__5411 (
            .O(N__22101),
            .I(N__22087));
    CascadeMux I__5410 (
            .O(N__22100),
            .I(N__22084));
    InMux I__5409 (
            .O(N__22097),
            .I(N__22081));
    InMux I__5408 (
            .O(N__22096),
            .I(N__22078));
    CascadeMux I__5407 (
            .O(N__22095),
            .I(N__22074));
    CascadeMux I__5406 (
            .O(N__22094),
            .I(N__22070));
    CascadeMux I__5405 (
            .O(N__22093),
            .I(N__22066));
    CascadeMux I__5404 (
            .O(N__22092),
            .I(N__22062));
    CascadeMux I__5403 (
            .O(N__22091),
            .I(N__22059));
    InMux I__5402 (
            .O(N__22090),
            .I(N__22056));
    InMux I__5401 (
            .O(N__22087),
            .I(N__22051));
    InMux I__5400 (
            .O(N__22084),
            .I(N__22051));
    LocalMux I__5399 (
            .O(N__22081),
            .I(N__22046));
    LocalMux I__5398 (
            .O(N__22078),
            .I(N__22046));
    InMux I__5397 (
            .O(N__22077),
            .I(N__22041));
    InMux I__5396 (
            .O(N__22074),
            .I(N__22041));
    InMux I__5395 (
            .O(N__22073),
            .I(N__22036));
    InMux I__5394 (
            .O(N__22070),
            .I(N__22036));
    CascadeMux I__5393 (
            .O(N__22069),
            .I(N__22033));
    InMux I__5392 (
            .O(N__22066),
            .I(N__22030));
    CascadeMux I__5391 (
            .O(N__22065),
            .I(N__22027));
    InMux I__5390 (
            .O(N__22062),
            .I(N__22024));
    InMux I__5389 (
            .O(N__22059),
            .I(N__22021));
    LocalMux I__5388 (
            .O(N__22056),
            .I(N__22014));
    LocalMux I__5387 (
            .O(N__22051),
            .I(N__22014));
    Span4Mux_v I__5386 (
            .O(N__22046),
            .I(N__22014));
    LocalMux I__5385 (
            .O(N__22041),
            .I(N__22009));
    LocalMux I__5384 (
            .O(N__22036),
            .I(N__22009));
    InMux I__5383 (
            .O(N__22033),
            .I(N__22006));
    LocalMux I__5382 (
            .O(N__22030),
            .I(N__22003));
    InMux I__5381 (
            .O(N__22027),
            .I(N__22000));
    LocalMux I__5380 (
            .O(N__22024),
            .I(N__21997));
    LocalMux I__5379 (
            .O(N__22021),
            .I(N__21990));
    Span4Mux_v I__5378 (
            .O(N__22014),
            .I(N__21990));
    Span4Mux_v I__5377 (
            .O(N__22009),
            .I(N__21990));
    LocalMux I__5376 (
            .O(N__22006),
            .I(N__21985));
    Span4Mux_h I__5375 (
            .O(N__22003),
            .I(N__21985));
    LocalMux I__5374 (
            .O(N__22000),
            .I(\Lab_UT.scctrl.state_i_3_0_rep2 ));
    Odrv12 I__5373 (
            .O(N__21997),
            .I(\Lab_UT.scctrl.state_i_3_0_rep2 ));
    Odrv4 I__5372 (
            .O(N__21990),
            .I(\Lab_UT.scctrl.state_i_3_0_rep2 ));
    Odrv4 I__5371 (
            .O(N__21985),
            .I(\Lab_UT.scctrl.state_i_3_0_rep2 ));
    InMux I__5370 (
            .O(N__21976),
            .I(N__21972));
    InMux I__5369 (
            .O(N__21975),
            .I(N__21969));
    LocalMux I__5368 (
            .O(N__21972),
            .I(N__21964));
    LocalMux I__5367 (
            .O(N__21969),
            .I(N__21964));
    Odrv4 I__5366 (
            .O(N__21964),
            .I(rst_i_3_fast));
    InMux I__5365 (
            .O(N__21961),
            .I(N__21958));
    LocalMux I__5364 (
            .O(N__21958),
            .I(\Lab_UT.scctrl.g1_i_0 ));
    InMux I__5363 (
            .O(N__21955),
            .I(N__21952));
    LocalMux I__5362 (
            .O(N__21952),
            .I(N__21944));
    InMux I__5361 (
            .O(N__21951),
            .I(N__21938));
    InMux I__5360 (
            .O(N__21950),
            .I(N__21933));
    InMux I__5359 (
            .O(N__21949),
            .I(N__21933));
    InMux I__5358 (
            .O(N__21948),
            .I(N__21930));
    InMux I__5357 (
            .O(N__21947),
            .I(N__21924));
    Span4Mux_s1_v I__5356 (
            .O(N__21944),
            .I(N__21919));
    InMux I__5355 (
            .O(N__21943),
            .I(N__21916));
    InMux I__5354 (
            .O(N__21942),
            .I(N__21913));
    InMux I__5353 (
            .O(N__21941),
            .I(N__21910));
    LocalMux I__5352 (
            .O(N__21938),
            .I(N__21907));
    LocalMux I__5351 (
            .O(N__21933),
            .I(N__21904));
    LocalMux I__5350 (
            .O(N__21930),
            .I(N__21901));
    InMux I__5349 (
            .O(N__21929),
            .I(N__21896));
    InMux I__5348 (
            .O(N__21928),
            .I(N__21896));
    InMux I__5347 (
            .O(N__21927),
            .I(N__21893));
    LocalMux I__5346 (
            .O(N__21924),
            .I(N__21890));
    InMux I__5345 (
            .O(N__21923),
            .I(N__21887));
    InMux I__5344 (
            .O(N__21922),
            .I(N__21884));
    Span4Mux_h I__5343 (
            .O(N__21919),
            .I(N__21879));
    LocalMux I__5342 (
            .O(N__21916),
            .I(N__21879));
    LocalMux I__5341 (
            .O(N__21913),
            .I(N__21874));
    LocalMux I__5340 (
            .O(N__21910),
            .I(N__21874));
    Span4Mux_v I__5339 (
            .O(N__21907),
            .I(N__21871));
    Span4Mux_h I__5338 (
            .O(N__21904),
            .I(N__21862));
    Span4Mux_s2_h I__5337 (
            .O(N__21901),
            .I(N__21862));
    LocalMux I__5336 (
            .O(N__21896),
            .I(N__21859));
    LocalMux I__5335 (
            .O(N__21893),
            .I(N__21856));
    Span12Mux_s11_h I__5334 (
            .O(N__21890),
            .I(N__21853));
    LocalMux I__5333 (
            .O(N__21887),
            .I(N__21850));
    LocalMux I__5332 (
            .O(N__21884),
            .I(N__21843));
    Span4Mux_v I__5331 (
            .O(N__21879),
            .I(N__21843));
    Span4Mux_h I__5330 (
            .O(N__21874),
            .I(N__21843));
    Span4Mux_v I__5329 (
            .O(N__21871),
            .I(N__21840));
    InMux I__5328 (
            .O(N__21870),
            .I(N__21837));
    InMux I__5327 (
            .O(N__21869),
            .I(N__21830));
    InMux I__5326 (
            .O(N__21868),
            .I(N__21830));
    InMux I__5325 (
            .O(N__21867),
            .I(N__21830));
    Span4Mux_v I__5324 (
            .O(N__21862),
            .I(N__21823));
    Span4Mux_s2_h I__5323 (
            .O(N__21859),
            .I(N__21823));
    Span4Mux_h I__5322 (
            .O(N__21856),
            .I(N__21823));
    Span12Mux_v I__5321 (
            .O(N__21853),
            .I(N__21820));
    Span4Mux_s2_h I__5320 (
            .O(N__21850),
            .I(N__21815));
    Span4Mux_v I__5319 (
            .O(N__21843),
            .I(N__21815));
    Odrv4 I__5318 (
            .O(N__21840),
            .I(\Lab_UT.state_i_3_0 ));
    LocalMux I__5317 (
            .O(N__21837),
            .I(\Lab_UT.state_i_3_0 ));
    LocalMux I__5316 (
            .O(N__21830),
            .I(\Lab_UT.state_i_3_0 ));
    Odrv4 I__5315 (
            .O(N__21823),
            .I(\Lab_UT.state_i_3_0 ));
    Odrv12 I__5314 (
            .O(N__21820),
            .I(\Lab_UT.state_i_3_0 ));
    Odrv4 I__5313 (
            .O(N__21815),
            .I(\Lab_UT.state_i_3_0 ));
    CascadeMux I__5312 (
            .O(N__21802),
            .I(N__21799));
    InMux I__5311 (
            .O(N__21799),
            .I(N__21796));
    LocalMux I__5310 (
            .O(N__21796),
            .I(\Lab_UT.scctrl.g0_0_i_a8_3_1 ));
    CascadeMux I__5309 (
            .O(N__21793),
            .I(N__21784));
    CascadeMux I__5308 (
            .O(N__21792),
            .I(N__21779));
    CascadeMux I__5307 (
            .O(N__21791),
            .I(N__21776));
    InMux I__5306 (
            .O(N__21790),
            .I(N__21771));
    InMux I__5305 (
            .O(N__21789),
            .I(N__21771));
    InMux I__5304 (
            .O(N__21788),
            .I(N__21757));
    InMux I__5303 (
            .O(N__21787),
            .I(N__21753));
    InMux I__5302 (
            .O(N__21784),
            .I(N__21750));
    InMux I__5301 (
            .O(N__21783),
            .I(N__21747));
    CascadeMux I__5300 (
            .O(N__21782),
            .I(N__21744));
    InMux I__5299 (
            .O(N__21779),
            .I(N__21739));
    InMux I__5298 (
            .O(N__21776),
            .I(N__21736));
    LocalMux I__5297 (
            .O(N__21771),
            .I(N__21732));
    InMux I__5296 (
            .O(N__21770),
            .I(N__21729));
    InMux I__5295 (
            .O(N__21769),
            .I(N__21726));
    InMux I__5294 (
            .O(N__21768),
            .I(N__21723));
    InMux I__5293 (
            .O(N__21767),
            .I(N__21716));
    InMux I__5292 (
            .O(N__21766),
            .I(N__21716));
    InMux I__5291 (
            .O(N__21765),
            .I(N__21716));
    InMux I__5290 (
            .O(N__21764),
            .I(N__21707));
    InMux I__5289 (
            .O(N__21763),
            .I(N__21707));
    InMux I__5288 (
            .O(N__21762),
            .I(N__21707));
    InMux I__5287 (
            .O(N__21761),
            .I(N__21702));
    InMux I__5286 (
            .O(N__21760),
            .I(N__21702));
    LocalMux I__5285 (
            .O(N__21757),
            .I(N__21699));
    InMux I__5284 (
            .O(N__21756),
            .I(N__21695));
    LocalMux I__5283 (
            .O(N__21753),
            .I(N__21692));
    LocalMux I__5282 (
            .O(N__21750),
            .I(N__21689));
    LocalMux I__5281 (
            .O(N__21747),
            .I(N__21685));
    InMux I__5280 (
            .O(N__21744),
            .I(N__21682));
    InMux I__5279 (
            .O(N__21743),
            .I(N__21677));
    InMux I__5278 (
            .O(N__21742),
            .I(N__21677));
    LocalMux I__5277 (
            .O(N__21739),
            .I(N__21674));
    LocalMux I__5276 (
            .O(N__21736),
            .I(N__21670));
    CascadeMux I__5275 (
            .O(N__21735),
            .I(N__21665));
    Span4Mux_v I__5274 (
            .O(N__21732),
            .I(N__21662));
    LocalMux I__5273 (
            .O(N__21729),
            .I(N__21659));
    LocalMux I__5272 (
            .O(N__21726),
            .I(N__21656));
    LocalMux I__5271 (
            .O(N__21723),
            .I(N__21651));
    LocalMux I__5270 (
            .O(N__21716),
            .I(N__21651));
    InMux I__5269 (
            .O(N__21715),
            .I(N__21646));
    InMux I__5268 (
            .O(N__21714),
            .I(N__21646));
    LocalMux I__5267 (
            .O(N__21707),
            .I(N__21641));
    LocalMux I__5266 (
            .O(N__21702),
            .I(N__21641));
    Span4Mux_h I__5265 (
            .O(N__21699),
            .I(N__21638));
    InMux I__5264 (
            .O(N__21698),
            .I(N__21635));
    LocalMux I__5263 (
            .O(N__21695),
            .I(N__21628));
    Span4Mux_v I__5262 (
            .O(N__21692),
            .I(N__21628));
    Span4Mux_s1_h I__5261 (
            .O(N__21689),
            .I(N__21628));
    InMux I__5260 (
            .O(N__21688),
            .I(N__21625));
    Span12Mux_s5_h I__5259 (
            .O(N__21685),
            .I(N__21618));
    LocalMux I__5258 (
            .O(N__21682),
            .I(N__21618));
    LocalMux I__5257 (
            .O(N__21677),
            .I(N__21618));
    Span4Mux_v I__5256 (
            .O(N__21674),
            .I(N__21615));
    InMux I__5255 (
            .O(N__21673),
            .I(N__21612));
    Span4Mux_v I__5254 (
            .O(N__21670),
            .I(N__21609));
    InMux I__5253 (
            .O(N__21669),
            .I(N__21602));
    InMux I__5252 (
            .O(N__21668),
            .I(N__21602));
    InMux I__5251 (
            .O(N__21665),
            .I(N__21602));
    Span4Mux_h I__5250 (
            .O(N__21662),
            .I(N__21593));
    Span4Mux_h I__5249 (
            .O(N__21659),
            .I(N__21593));
    Span4Mux_h I__5248 (
            .O(N__21656),
            .I(N__21593));
    Span4Mux_v I__5247 (
            .O(N__21651),
            .I(N__21593));
    LocalMux I__5246 (
            .O(N__21646),
            .I(N__21588));
    Span4Mux_v I__5245 (
            .O(N__21641),
            .I(N__21588));
    Span4Mux_v I__5244 (
            .O(N__21638),
            .I(N__21581));
    LocalMux I__5243 (
            .O(N__21635),
            .I(N__21581));
    Span4Mux_h I__5242 (
            .O(N__21628),
            .I(N__21581));
    LocalMux I__5241 (
            .O(N__21625),
            .I(\Lab_UT.state_1 ));
    Odrv12 I__5240 (
            .O(N__21618),
            .I(\Lab_UT.state_1 ));
    Odrv4 I__5239 (
            .O(N__21615),
            .I(\Lab_UT.state_1 ));
    LocalMux I__5238 (
            .O(N__21612),
            .I(\Lab_UT.state_1 ));
    Odrv4 I__5237 (
            .O(N__21609),
            .I(\Lab_UT.state_1 ));
    LocalMux I__5236 (
            .O(N__21602),
            .I(\Lab_UT.state_1 ));
    Odrv4 I__5235 (
            .O(N__21593),
            .I(\Lab_UT.state_1 ));
    Odrv4 I__5234 (
            .O(N__21588),
            .I(\Lab_UT.state_1 ));
    Odrv4 I__5233 (
            .O(N__21581),
            .I(\Lab_UT.state_1 ));
    InMux I__5232 (
            .O(N__21562),
            .I(N__21559));
    LocalMux I__5231 (
            .O(N__21559),
            .I(\Lab_UT.scctrl.state_1_RNO_3Z0Z_0 ));
    InMux I__5230 (
            .O(N__21556),
            .I(N__21553));
    LocalMux I__5229 (
            .O(N__21553),
            .I(N__21550));
    Odrv4 I__5228 (
            .O(N__21550),
            .I(\Lab_UT.scctrl.N_13_0 ));
    InMux I__5227 (
            .O(N__21547),
            .I(N__21543));
    InMux I__5226 (
            .O(N__21546),
            .I(N__21540));
    LocalMux I__5225 (
            .O(N__21543),
            .I(N__21537));
    LocalMux I__5224 (
            .O(N__21540),
            .I(N__21534));
    Span4Mux_s0_h I__5223 (
            .O(N__21537),
            .I(N__21531));
    Span4Mux_h I__5222 (
            .O(N__21534),
            .I(N__21525));
    Span4Mux_h I__5221 (
            .O(N__21531),
            .I(N__21522));
    InMux I__5220 (
            .O(N__21530),
            .I(N__21515));
    InMux I__5219 (
            .O(N__21529),
            .I(N__21515));
    InMux I__5218 (
            .O(N__21528),
            .I(N__21515));
    Odrv4 I__5217 (
            .O(N__21525),
            .I(\Lab_UT.N_191 ));
    Odrv4 I__5216 (
            .O(N__21522),
            .I(\Lab_UT.N_191 ));
    LocalMux I__5215 (
            .O(N__21515),
            .I(\Lab_UT.N_191 ));
    CascadeMux I__5214 (
            .O(N__21508),
            .I(N__21505));
    InMux I__5213 (
            .O(N__21505),
            .I(N__21502));
    LocalMux I__5212 (
            .O(N__21502),
            .I(N__21499));
    Span4Mux_s1_h I__5211 (
            .O(N__21499),
            .I(N__21496));
    Span4Mux_h I__5210 (
            .O(N__21496),
            .I(N__21493));
    Odrv4 I__5209 (
            .O(N__21493),
            .I(\Lab_UT.scctrl.G_24_i_a4_0_1 ));
    InMux I__5208 (
            .O(N__21490),
            .I(N__21486));
    InMux I__5207 (
            .O(N__21489),
            .I(N__21483));
    LocalMux I__5206 (
            .O(N__21486),
            .I(N__21480));
    LocalMux I__5205 (
            .O(N__21483),
            .I(N__21474));
    Span4Mux_v I__5204 (
            .O(N__21480),
            .I(N__21471));
    InMux I__5203 (
            .O(N__21479),
            .I(N__21464));
    InMux I__5202 (
            .O(N__21478),
            .I(N__21464));
    InMux I__5201 (
            .O(N__21477),
            .I(N__21464));
    Span4Mux_h I__5200 (
            .O(N__21474),
            .I(N__21457));
    Span4Mux_h I__5199 (
            .O(N__21471),
            .I(N__21457));
    LocalMux I__5198 (
            .O(N__21464),
            .I(N__21457));
    Odrv4 I__5197 (
            .O(N__21457),
            .I(\Lab_UT.next_state_1_0_0_3 ));
    InMux I__5196 (
            .O(N__21454),
            .I(N__21451));
    LocalMux I__5195 (
            .O(N__21451),
            .I(N__21448));
    Odrv4 I__5194 (
            .O(N__21448),
            .I(\Lab_UT.scctrl.N_10_2 ));
    InMux I__5193 (
            .O(N__21445),
            .I(N__21441));
    CascadeMux I__5192 (
            .O(N__21444),
            .I(N__21436));
    LocalMux I__5191 (
            .O(N__21441),
            .I(N__21433));
    CascadeMux I__5190 (
            .O(N__21440),
            .I(N__21429));
    CascadeMux I__5189 (
            .O(N__21439),
            .I(N__21421));
    InMux I__5188 (
            .O(N__21436),
            .I(N__21416));
    Span4Mux_v I__5187 (
            .O(N__21433),
            .I(N__21413));
    InMux I__5186 (
            .O(N__21432),
            .I(N__21410));
    InMux I__5185 (
            .O(N__21429),
            .I(N__21402));
    InMux I__5184 (
            .O(N__21428),
            .I(N__21402));
    InMux I__5183 (
            .O(N__21427),
            .I(N__21392));
    InMux I__5182 (
            .O(N__21426),
            .I(N__21392));
    CascadeMux I__5181 (
            .O(N__21425),
            .I(N__21389));
    InMux I__5180 (
            .O(N__21424),
            .I(N__21383));
    InMux I__5179 (
            .O(N__21421),
            .I(N__21383));
    InMux I__5178 (
            .O(N__21420),
            .I(N__21378));
    InMux I__5177 (
            .O(N__21419),
            .I(N__21378));
    LocalMux I__5176 (
            .O(N__21416),
            .I(N__21369));
    Span4Mux_v I__5175 (
            .O(N__21413),
            .I(N__21369));
    LocalMux I__5174 (
            .O(N__21410),
            .I(N__21369));
    InMux I__5173 (
            .O(N__21409),
            .I(N__21364));
    InMux I__5172 (
            .O(N__21408),
            .I(N__21364));
    InMux I__5171 (
            .O(N__21407),
            .I(N__21359));
    LocalMux I__5170 (
            .O(N__21402),
            .I(N__21356));
    InMux I__5169 (
            .O(N__21401),
            .I(N__21351));
    InMux I__5168 (
            .O(N__21400),
            .I(N__21351));
    InMux I__5167 (
            .O(N__21399),
            .I(N__21344));
    InMux I__5166 (
            .O(N__21398),
            .I(N__21344));
    InMux I__5165 (
            .O(N__21397),
            .I(N__21344));
    LocalMux I__5164 (
            .O(N__21392),
            .I(N__21341));
    InMux I__5163 (
            .O(N__21389),
            .I(N__21336));
    InMux I__5162 (
            .O(N__21388),
            .I(N__21336));
    LocalMux I__5161 (
            .O(N__21383),
            .I(N__21331));
    LocalMux I__5160 (
            .O(N__21378),
            .I(N__21331));
    InMux I__5159 (
            .O(N__21377),
            .I(N__21328));
    InMux I__5158 (
            .O(N__21376),
            .I(N__21325));
    Span4Mux_v I__5157 (
            .O(N__21369),
            .I(N__21321));
    LocalMux I__5156 (
            .O(N__21364),
            .I(N__21318));
    InMux I__5155 (
            .O(N__21363),
            .I(N__21313));
    InMux I__5154 (
            .O(N__21362),
            .I(N__21313));
    LocalMux I__5153 (
            .O(N__21359),
            .I(N__21306));
    Span4Mux_h I__5152 (
            .O(N__21356),
            .I(N__21306));
    LocalMux I__5151 (
            .O(N__21351),
            .I(N__21306));
    LocalMux I__5150 (
            .O(N__21344),
            .I(N__21303));
    Span4Mux_v I__5149 (
            .O(N__21341),
            .I(N__21300));
    LocalMux I__5148 (
            .O(N__21336),
            .I(N__21291));
    Span4Mux_v I__5147 (
            .O(N__21331),
            .I(N__21291));
    LocalMux I__5146 (
            .O(N__21328),
            .I(N__21291));
    LocalMux I__5145 (
            .O(N__21325),
            .I(N__21291));
    InMux I__5144 (
            .O(N__21324),
            .I(N__21287));
    Span4Mux_v I__5143 (
            .O(N__21321),
            .I(N__21284));
    Span4Mux_h I__5142 (
            .O(N__21318),
            .I(N__21277));
    LocalMux I__5141 (
            .O(N__21313),
            .I(N__21277));
    Span4Mux_h I__5140 (
            .O(N__21306),
            .I(N__21277));
    Span4Mux_h I__5139 (
            .O(N__21303),
            .I(N__21272));
    Span4Mux_h I__5138 (
            .O(N__21300),
            .I(N__21272));
    Span4Mux_h I__5137 (
            .O(N__21291),
            .I(N__21269));
    InMux I__5136 (
            .O(N__21290),
            .I(N__21266));
    LocalMux I__5135 (
            .O(N__21287),
            .I(\Lab_UT.N_169_0 ));
    Odrv4 I__5134 (
            .O(N__21284),
            .I(\Lab_UT.N_169_0 ));
    Odrv4 I__5133 (
            .O(N__21277),
            .I(\Lab_UT.N_169_0 ));
    Odrv4 I__5132 (
            .O(N__21272),
            .I(\Lab_UT.N_169_0 ));
    Odrv4 I__5131 (
            .O(N__21269),
            .I(\Lab_UT.N_169_0 ));
    LocalMux I__5130 (
            .O(N__21266),
            .I(\Lab_UT.N_169_0 ));
    InMux I__5129 (
            .O(N__21253),
            .I(N__21250));
    LocalMux I__5128 (
            .O(N__21250),
            .I(N__21245));
    InMux I__5127 (
            .O(N__21249),
            .I(N__21242));
    InMux I__5126 (
            .O(N__21248),
            .I(N__21239));
    Span4Mux_v I__5125 (
            .O(N__21245),
            .I(N__21236));
    LocalMux I__5124 (
            .O(N__21242),
            .I(N__21233));
    LocalMux I__5123 (
            .O(N__21239),
            .I(N__21230));
    Span4Mux_v I__5122 (
            .O(N__21236),
            .I(N__21227));
    Span12Mux_v I__5121 (
            .O(N__21233),
            .I(N__21224));
    Span4Mux_h I__5120 (
            .O(N__21230),
            .I(N__21221));
    Odrv4 I__5119 (
            .O(N__21227),
            .I(\Lab_UT.scctrl.N_223_1 ));
    Odrv12 I__5118 (
            .O(N__21224),
            .I(\Lab_UT.scctrl.N_223_1 ));
    Odrv4 I__5117 (
            .O(N__21221),
            .I(\Lab_UT.scctrl.N_223_1 ));
    IoInMux I__5116 (
            .O(N__21214),
            .I(N__21211));
    LocalMux I__5115 (
            .O(N__21211),
            .I(led_c_4));
    CascadeMux I__5114 (
            .O(N__21208),
            .I(N__21203));
    CascadeMux I__5113 (
            .O(N__21207),
            .I(N__21197));
    InMux I__5112 (
            .O(N__21206),
            .I(N__21192));
    InMux I__5111 (
            .O(N__21203),
            .I(N__21186));
    CascadeMux I__5110 (
            .O(N__21202),
            .I(N__21182));
    CascadeMux I__5109 (
            .O(N__21201),
            .I(N__21179));
    CascadeMux I__5108 (
            .O(N__21200),
            .I(N__21176));
    InMux I__5107 (
            .O(N__21197),
            .I(N__21169));
    InMux I__5106 (
            .O(N__21196),
            .I(N__21166));
    CascadeMux I__5105 (
            .O(N__21195),
            .I(N__21162));
    LocalMux I__5104 (
            .O(N__21192),
            .I(N__21157));
    InMux I__5103 (
            .O(N__21191),
            .I(N__21152));
    InMux I__5102 (
            .O(N__21190),
            .I(N__21152));
    InMux I__5101 (
            .O(N__21189),
            .I(N__21149));
    LocalMux I__5100 (
            .O(N__21186),
            .I(N__21146));
    InMux I__5099 (
            .O(N__21185),
            .I(N__21143));
    InMux I__5098 (
            .O(N__21182),
            .I(N__21138));
    InMux I__5097 (
            .O(N__21179),
            .I(N__21138));
    InMux I__5096 (
            .O(N__21176),
            .I(N__21135));
    InMux I__5095 (
            .O(N__21175),
            .I(N__21130));
    InMux I__5094 (
            .O(N__21174),
            .I(N__21130));
    CascadeMux I__5093 (
            .O(N__21173),
            .I(N__21123));
    CascadeMux I__5092 (
            .O(N__21172),
            .I(N__21120));
    LocalMux I__5091 (
            .O(N__21169),
            .I(N__21117));
    LocalMux I__5090 (
            .O(N__21166),
            .I(N__21114));
    InMux I__5089 (
            .O(N__21165),
            .I(N__21109));
    InMux I__5088 (
            .O(N__21162),
            .I(N__21109));
    InMux I__5087 (
            .O(N__21161),
            .I(N__21104));
    InMux I__5086 (
            .O(N__21160),
            .I(N__21104));
    Span4Mux_s3_h I__5085 (
            .O(N__21157),
            .I(N__21095));
    LocalMux I__5084 (
            .O(N__21152),
            .I(N__21095));
    LocalMux I__5083 (
            .O(N__21149),
            .I(N__21095));
    Span4Mux_h I__5082 (
            .O(N__21146),
            .I(N__21095));
    LocalMux I__5081 (
            .O(N__21143),
            .I(N__21092));
    LocalMux I__5080 (
            .O(N__21138),
            .I(N__21087));
    LocalMux I__5079 (
            .O(N__21135),
            .I(N__21087));
    LocalMux I__5078 (
            .O(N__21130),
            .I(N__21084));
    CascadeMux I__5077 (
            .O(N__21129),
            .I(N__21081));
    CascadeMux I__5076 (
            .O(N__21128),
            .I(N__21078));
    InMux I__5075 (
            .O(N__21127),
            .I(N__21075));
    InMux I__5074 (
            .O(N__21126),
            .I(N__21072));
    InMux I__5073 (
            .O(N__21123),
            .I(N__21069));
    InMux I__5072 (
            .O(N__21120),
            .I(N__21066));
    Span12Mux_s4_h I__5071 (
            .O(N__21117),
            .I(N__21059));
    Span12Mux_s8_v I__5070 (
            .O(N__21114),
            .I(N__21059));
    LocalMux I__5069 (
            .O(N__21109),
            .I(N__21059));
    LocalMux I__5068 (
            .O(N__21104),
            .I(N__21054));
    Span4Mux_v I__5067 (
            .O(N__21095),
            .I(N__21054));
    Span4Mux_v I__5066 (
            .O(N__21092),
            .I(N__21047));
    Span4Mux_v I__5065 (
            .O(N__21087),
            .I(N__21047));
    Span4Mux_v I__5064 (
            .O(N__21084),
            .I(N__21047));
    InMux I__5063 (
            .O(N__21081),
            .I(N__21042));
    InMux I__5062 (
            .O(N__21078),
            .I(N__21042));
    LocalMux I__5061 (
            .O(N__21075),
            .I(\Lab_UT.un1_state_3_1 ));
    LocalMux I__5060 (
            .O(N__21072),
            .I(\Lab_UT.un1_state_3_1 ));
    LocalMux I__5059 (
            .O(N__21069),
            .I(\Lab_UT.un1_state_3_1 ));
    LocalMux I__5058 (
            .O(N__21066),
            .I(\Lab_UT.un1_state_3_1 ));
    Odrv12 I__5057 (
            .O(N__21059),
            .I(\Lab_UT.un1_state_3_1 ));
    Odrv4 I__5056 (
            .O(N__21054),
            .I(\Lab_UT.un1_state_3_1 ));
    Odrv4 I__5055 (
            .O(N__21047),
            .I(\Lab_UT.un1_state_3_1 ));
    LocalMux I__5054 (
            .O(N__21042),
            .I(\Lab_UT.un1_state_3_1 ));
    InMux I__5053 (
            .O(N__21025),
            .I(N__21016));
    InMux I__5052 (
            .O(N__21024),
            .I(N__21008));
    InMux I__5051 (
            .O(N__21023),
            .I(N__21003));
    InMux I__5050 (
            .O(N__21022),
            .I(N__21000));
    InMux I__5049 (
            .O(N__21021),
            .I(N__20997));
    InMux I__5048 (
            .O(N__21020),
            .I(N__20992));
    InMux I__5047 (
            .O(N__21019),
            .I(N__20992));
    LocalMux I__5046 (
            .O(N__21016),
            .I(N__20978));
    InMux I__5045 (
            .O(N__21015),
            .I(N__20975));
    InMux I__5044 (
            .O(N__21014),
            .I(N__20972));
    CascadeMux I__5043 (
            .O(N__21013),
            .I(N__20969));
    InMux I__5042 (
            .O(N__21012),
            .I(N__20964));
    InMux I__5041 (
            .O(N__21011),
            .I(N__20964));
    LocalMux I__5040 (
            .O(N__21008),
            .I(N__20961));
    InMux I__5039 (
            .O(N__21007),
            .I(N__20956));
    InMux I__5038 (
            .O(N__21006),
            .I(N__20956));
    LocalMux I__5037 (
            .O(N__21003),
            .I(N__20953));
    LocalMux I__5036 (
            .O(N__21000),
            .I(N__20948));
    LocalMux I__5035 (
            .O(N__20997),
            .I(N__20948));
    LocalMux I__5034 (
            .O(N__20992),
            .I(N__20945));
    InMux I__5033 (
            .O(N__20991),
            .I(N__20940));
    InMux I__5032 (
            .O(N__20990),
            .I(N__20940));
    InMux I__5031 (
            .O(N__20989),
            .I(N__20937));
    InMux I__5030 (
            .O(N__20988),
            .I(N__20932));
    InMux I__5029 (
            .O(N__20987),
            .I(N__20932));
    InMux I__5028 (
            .O(N__20986),
            .I(N__20920));
    InMux I__5027 (
            .O(N__20985),
            .I(N__20920));
    InMux I__5026 (
            .O(N__20984),
            .I(N__20920));
    InMux I__5025 (
            .O(N__20983),
            .I(N__20913));
    InMux I__5024 (
            .O(N__20982),
            .I(N__20913));
    InMux I__5023 (
            .O(N__20981),
            .I(N__20913));
    Span4Mux_s1_h I__5022 (
            .O(N__20978),
            .I(N__20905));
    LocalMux I__5021 (
            .O(N__20975),
            .I(N__20905));
    LocalMux I__5020 (
            .O(N__20972),
            .I(N__20902));
    InMux I__5019 (
            .O(N__20969),
            .I(N__20899));
    LocalMux I__5018 (
            .O(N__20964),
            .I(N__20892));
    Span4Mux_h I__5017 (
            .O(N__20961),
            .I(N__20892));
    LocalMux I__5016 (
            .O(N__20956),
            .I(N__20892));
    Span4Mux_v I__5015 (
            .O(N__20953),
            .I(N__20883));
    Span4Mux_v I__5014 (
            .O(N__20948),
            .I(N__20883));
    Span4Mux_h I__5013 (
            .O(N__20945),
            .I(N__20883));
    LocalMux I__5012 (
            .O(N__20940),
            .I(N__20883));
    LocalMux I__5011 (
            .O(N__20937),
            .I(N__20878));
    LocalMux I__5010 (
            .O(N__20932),
            .I(N__20878));
    InMux I__5009 (
            .O(N__20931),
            .I(N__20871));
    InMux I__5008 (
            .O(N__20930),
            .I(N__20871));
    InMux I__5007 (
            .O(N__20929),
            .I(N__20871));
    InMux I__5006 (
            .O(N__20928),
            .I(N__20866));
    InMux I__5005 (
            .O(N__20927),
            .I(N__20866));
    LocalMux I__5004 (
            .O(N__20920),
            .I(N__20861));
    LocalMux I__5003 (
            .O(N__20913),
            .I(N__20861));
    InMux I__5002 (
            .O(N__20912),
            .I(N__20854));
    InMux I__5001 (
            .O(N__20911),
            .I(N__20854));
    InMux I__5000 (
            .O(N__20910),
            .I(N__20854));
    Span4Mux_h I__4999 (
            .O(N__20905),
            .I(N__20847));
    Span4Mux_v I__4998 (
            .O(N__20902),
            .I(N__20847));
    LocalMux I__4997 (
            .O(N__20899),
            .I(N__20847));
    Odrv4 I__4996 (
            .O(N__20892),
            .I(L4_PrintBuf));
    Odrv4 I__4995 (
            .O(N__20883),
            .I(L4_PrintBuf));
    Odrv4 I__4994 (
            .O(N__20878),
            .I(L4_PrintBuf));
    LocalMux I__4993 (
            .O(N__20871),
            .I(L4_PrintBuf));
    LocalMux I__4992 (
            .O(N__20866),
            .I(L4_PrintBuf));
    Odrv12 I__4991 (
            .O(N__20861),
            .I(L4_PrintBuf));
    LocalMux I__4990 (
            .O(N__20854),
            .I(L4_PrintBuf));
    Odrv4 I__4989 (
            .O(N__20847),
            .I(L4_PrintBuf));
    InMux I__4988 (
            .O(N__20830),
            .I(N__20827));
    LocalMux I__4987 (
            .O(N__20827),
            .I(N__20824));
    Span4Mux_h I__4986 (
            .O(N__20824),
            .I(N__20821));
    Odrv4 I__4985 (
            .O(N__20821),
            .I(\Lab_UT.scctrl.m26_i_o4_1_2 ));
    CascadeMux I__4984 (
            .O(N__20818),
            .I(\Lab_UT.scctrl.G_24_i_o3_0_0_cascade_ ));
    CascadeMux I__4983 (
            .O(N__20815),
            .I(N__20811));
    InMux I__4982 (
            .O(N__20814),
            .I(N__20800));
    InMux I__4981 (
            .O(N__20811),
            .I(N__20797));
    InMux I__4980 (
            .O(N__20810),
            .I(N__20792));
    InMux I__4979 (
            .O(N__20809),
            .I(N__20792));
    InMux I__4978 (
            .O(N__20808),
            .I(N__20788));
    InMux I__4977 (
            .O(N__20807),
            .I(N__20781));
    InMux I__4976 (
            .O(N__20806),
            .I(N__20776));
    InMux I__4975 (
            .O(N__20805),
            .I(N__20776));
    InMux I__4974 (
            .O(N__20804),
            .I(N__20771));
    InMux I__4973 (
            .O(N__20803),
            .I(N__20771));
    LocalMux I__4972 (
            .O(N__20800),
            .I(N__20768));
    LocalMux I__4971 (
            .O(N__20797),
            .I(N__20765));
    LocalMux I__4970 (
            .O(N__20792),
            .I(N__20762));
    InMux I__4969 (
            .O(N__20791),
            .I(N__20759));
    LocalMux I__4968 (
            .O(N__20788),
            .I(N__20754));
    InMux I__4967 (
            .O(N__20787),
            .I(N__20749));
    InMux I__4966 (
            .O(N__20786),
            .I(N__20742));
    InMux I__4965 (
            .O(N__20785),
            .I(N__20742));
    InMux I__4964 (
            .O(N__20784),
            .I(N__20742));
    LocalMux I__4963 (
            .O(N__20781),
            .I(N__20737));
    LocalMux I__4962 (
            .O(N__20776),
            .I(N__20737));
    LocalMux I__4961 (
            .O(N__20771),
            .I(N__20734));
    Span4Mux_s1_h I__4960 (
            .O(N__20768),
            .I(N__20729));
    Span4Mux_v I__4959 (
            .O(N__20765),
            .I(N__20729));
    Span4Mux_v I__4958 (
            .O(N__20762),
            .I(N__20726));
    LocalMux I__4957 (
            .O(N__20759),
            .I(N__20723));
    InMux I__4956 (
            .O(N__20758),
            .I(N__20720));
    CascadeMux I__4955 (
            .O(N__20757),
            .I(N__20714));
    Span4Mux_v I__4954 (
            .O(N__20754),
            .I(N__20710));
    InMux I__4953 (
            .O(N__20753),
            .I(N__20707));
    InMux I__4952 (
            .O(N__20752),
            .I(N__20704));
    LocalMux I__4951 (
            .O(N__20749),
            .I(N__20697));
    LocalMux I__4950 (
            .O(N__20742),
            .I(N__20697));
    Span4Mux_h I__4949 (
            .O(N__20737),
            .I(N__20697));
    Span4Mux_v I__4948 (
            .O(N__20734),
            .I(N__20692));
    Span4Mux_h I__4947 (
            .O(N__20729),
            .I(N__20692));
    Span4Mux_h I__4946 (
            .O(N__20726),
            .I(N__20685));
    Span4Mux_v I__4945 (
            .O(N__20723),
            .I(N__20685));
    LocalMux I__4944 (
            .O(N__20720),
            .I(N__20685));
    InMux I__4943 (
            .O(N__20719),
            .I(N__20682));
    InMux I__4942 (
            .O(N__20718),
            .I(N__20679));
    InMux I__4941 (
            .O(N__20717),
            .I(N__20676));
    InMux I__4940 (
            .O(N__20714),
            .I(N__20671));
    InMux I__4939 (
            .O(N__20713),
            .I(N__20671));
    Odrv4 I__4938 (
            .O(N__20710),
            .I(bu_rx_data_rdy));
    LocalMux I__4937 (
            .O(N__20707),
            .I(bu_rx_data_rdy));
    LocalMux I__4936 (
            .O(N__20704),
            .I(bu_rx_data_rdy));
    Odrv4 I__4935 (
            .O(N__20697),
            .I(bu_rx_data_rdy));
    Odrv4 I__4934 (
            .O(N__20692),
            .I(bu_rx_data_rdy));
    Odrv4 I__4933 (
            .O(N__20685),
            .I(bu_rx_data_rdy));
    LocalMux I__4932 (
            .O(N__20682),
            .I(bu_rx_data_rdy));
    LocalMux I__4931 (
            .O(N__20679),
            .I(bu_rx_data_rdy));
    LocalMux I__4930 (
            .O(N__20676),
            .I(bu_rx_data_rdy));
    LocalMux I__4929 (
            .O(N__20671),
            .I(bu_rx_data_rdy));
    CascadeMux I__4928 (
            .O(N__20650),
            .I(\Lab_UT.scctrl.N_6_5_cascade_ ));
    InMux I__4927 (
            .O(N__20647),
            .I(N__20644));
    LocalMux I__4926 (
            .O(N__20644),
            .I(\Lab_UT.scctrl.N_5_2 ));
    InMux I__4925 (
            .O(N__20641),
            .I(N__20638));
    LocalMux I__4924 (
            .O(N__20638),
            .I(N__20635));
    Odrv4 I__4923 (
            .O(N__20635),
            .I(\Lab_UT.scctrl.N_8_4 ));
    InMux I__4922 (
            .O(N__20632),
            .I(N__20627));
    InMux I__4921 (
            .O(N__20631),
            .I(N__20624));
    InMux I__4920 (
            .O(N__20630),
            .I(N__20621));
    LocalMux I__4919 (
            .O(N__20627),
            .I(N__20618));
    LocalMux I__4918 (
            .O(N__20624),
            .I(N__20615));
    LocalMux I__4917 (
            .O(N__20621),
            .I(N__20612));
    Span4Mux_h I__4916 (
            .O(N__20618),
            .I(N__20608));
    Span4Mux_v I__4915 (
            .O(N__20615),
            .I(N__20603));
    Span4Mux_v I__4914 (
            .O(N__20612),
            .I(N__20603));
    InMux I__4913 (
            .O(N__20611),
            .I(N__20600));
    Odrv4 I__4912 (
            .O(N__20608),
            .I(\Lab_UT.scctrl.N_4ctr ));
    Odrv4 I__4911 (
            .O(N__20603),
            .I(\Lab_UT.scctrl.N_4ctr ));
    LocalMux I__4910 (
            .O(N__20600),
            .I(\Lab_UT.scctrl.N_4ctr ));
    InMux I__4909 (
            .O(N__20593),
            .I(N__20590));
    LocalMux I__4908 (
            .O(N__20590),
            .I(N__20587));
    Span4Mux_h I__4907 (
            .O(N__20587),
            .I(N__20584));
    Span4Mux_v I__4906 (
            .O(N__20584),
            .I(N__20581));
    Odrv4 I__4905 (
            .O(N__20581),
            .I(\Lab_UT.scctrl.G_23_0_a9_1 ));
    InMux I__4904 (
            .O(N__20578),
            .I(N__20566));
    InMux I__4903 (
            .O(N__20577),
            .I(N__20557));
    InMux I__4902 (
            .O(N__20576),
            .I(N__20557));
    InMux I__4901 (
            .O(N__20575),
            .I(N__20551));
    InMux I__4900 (
            .O(N__20574),
            .I(N__20544));
    InMux I__4899 (
            .O(N__20573),
            .I(N__20544));
    InMux I__4898 (
            .O(N__20572),
            .I(N__20544));
    CascadeMux I__4897 (
            .O(N__20571),
            .I(N__20541));
    InMux I__4896 (
            .O(N__20570),
            .I(N__20532));
    InMux I__4895 (
            .O(N__20569),
            .I(N__20532));
    LocalMux I__4894 (
            .O(N__20566),
            .I(N__20527));
    InMux I__4893 (
            .O(N__20565),
            .I(N__20522));
    InMux I__4892 (
            .O(N__20564),
            .I(N__20522));
    InMux I__4891 (
            .O(N__20563),
            .I(N__20516));
    InMux I__4890 (
            .O(N__20562),
            .I(N__20516));
    LocalMux I__4889 (
            .O(N__20557),
            .I(N__20513));
    InMux I__4888 (
            .O(N__20556),
            .I(N__20505));
    InMux I__4887 (
            .O(N__20555),
            .I(N__20505));
    InMux I__4886 (
            .O(N__20554),
            .I(N__20505));
    LocalMux I__4885 (
            .O(N__20551),
            .I(N__20502));
    LocalMux I__4884 (
            .O(N__20544),
            .I(N__20499));
    InMux I__4883 (
            .O(N__20541),
            .I(N__20492));
    InMux I__4882 (
            .O(N__20540),
            .I(N__20492));
    InMux I__4881 (
            .O(N__20539),
            .I(N__20492));
    InMux I__4880 (
            .O(N__20538),
            .I(N__20489));
    InMux I__4879 (
            .O(N__20537),
            .I(N__20484));
    LocalMux I__4878 (
            .O(N__20532),
            .I(N__20481));
    InMux I__4877 (
            .O(N__20531),
            .I(N__20478));
    InMux I__4876 (
            .O(N__20530),
            .I(N__20475));
    Span4Mux_v I__4875 (
            .O(N__20527),
            .I(N__20470));
    LocalMux I__4874 (
            .O(N__20522),
            .I(N__20470));
    InMux I__4873 (
            .O(N__20521),
            .I(N__20467));
    LocalMux I__4872 (
            .O(N__20516),
            .I(N__20464));
    Span12Mux_s10_h I__4871 (
            .O(N__20513),
            .I(N__20459));
    CascadeMux I__4870 (
            .O(N__20512),
            .I(N__20455));
    LocalMux I__4869 (
            .O(N__20505),
            .I(N__20451));
    Span4Mux_s3_h I__4868 (
            .O(N__20502),
            .I(N__20444));
    Span4Mux_v I__4867 (
            .O(N__20499),
            .I(N__20444));
    LocalMux I__4866 (
            .O(N__20492),
            .I(N__20444));
    LocalMux I__4865 (
            .O(N__20489),
            .I(N__20439));
    InMux I__4864 (
            .O(N__20488),
            .I(N__20436));
    InMux I__4863 (
            .O(N__20487),
            .I(N__20433));
    LocalMux I__4862 (
            .O(N__20484),
            .I(N__20418));
    Span4Mux_h I__4861 (
            .O(N__20481),
            .I(N__20418));
    LocalMux I__4860 (
            .O(N__20478),
            .I(N__20418));
    LocalMux I__4859 (
            .O(N__20475),
            .I(N__20418));
    Span4Mux_h I__4858 (
            .O(N__20470),
            .I(N__20418));
    LocalMux I__4857 (
            .O(N__20467),
            .I(N__20418));
    Span4Mux_h I__4856 (
            .O(N__20464),
            .I(N__20418));
    InMux I__4855 (
            .O(N__20463),
            .I(N__20415));
    InMux I__4854 (
            .O(N__20462),
            .I(N__20412));
    Span12Mux_v I__4853 (
            .O(N__20459),
            .I(N__20409));
    InMux I__4852 (
            .O(N__20458),
            .I(N__20404));
    InMux I__4851 (
            .O(N__20455),
            .I(N__20404));
    InMux I__4850 (
            .O(N__20454),
            .I(N__20401));
    Span4Mux_s3_h I__4849 (
            .O(N__20451),
            .I(N__20396));
    Span4Mux_v I__4848 (
            .O(N__20444),
            .I(N__20396));
    InMux I__4847 (
            .O(N__20443),
            .I(N__20391));
    InMux I__4846 (
            .O(N__20442),
            .I(N__20391));
    Span12Mux_s2_v I__4845 (
            .O(N__20439),
            .I(N__20382));
    LocalMux I__4844 (
            .O(N__20436),
            .I(N__20382));
    LocalMux I__4843 (
            .O(N__20433),
            .I(N__20382));
    Sp12to4 I__4842 (
            .O(N__20418),
            .I(N__20382));
    LocalMux I__4841 (
            .O(N__20415),
            .I(\Lab_UT.state_i_3_1 ));
    LocalMux I__4840 (
            .O(N__20412),
            .I(\Lab_UT.state_i_3_1 ));
    Odrv12 I__4839 (
            .O(N__20409),
            .I(\Lab_UT.state_i_3_1 ));
    LocalMux I__4838 (
            .O(N__20404),
            .I(\Lab_UT.state_i_3_1 ));
    LocalMux I__4837 (
            .O(N__20401),
            .I(\Lab_UT.state_i_3_1 ));
    Odrv4 I__4836 (
            .O(N__20396),
            .I(\Lab_UT.state_i_3_1 ));
    LocalMux I__4835 (
            .O(N__20391),
            .I(\Lab_UT.state_i_3_1 ));
    Odrv12 I__4834 (
            .O(N__20382),
            .I(\Lab_UT.state_i_3_1 ));
    InMux I__4833 (
            .O(N__20365),
            .I(N__20356));
    InMux I__4832 (
            .O(N__20364),
            .I(N__20356));
    InMux I__4831 (
            .O(N__20363),
            .I(N__20356));
    LocalMux I__4830 (
            .O(N__20356),
            .I(N__20353));
    Odrv4 I__4829 (
            .O(N__20353),
            .I(\Lab_UT.scctrl.g0_i_a8_4_1 ));
    InMux I__4828 (
            .O(N__20350),
            .I(N__20345));
    CascadeMux I__4827 (
            .O(N__20349),
            .I(N__20342));
    InMux I__4826 (
            .O(N__20348),
            .I(N__20338));
    LocalMux I__4825 (
            .O(N__20345),
            .I(N__20335));
    InMux I__4824 (
            .O(N__20342),
            .I(N__20332));
    InMux I__4823 (
            .O(N__20341),
            .I(N__20328));
    LocalMux I__4822 (
            .O(N__20338),
            .I(N__20325));
    Span4Mux_s2_h I__4821 (
            .O(N__20335),
            .I(N__20320));
    LocalMux I__4820 (
            .O(N__20332),
            .I(N__20320));
    InMux I__4819 (
            .O(N__20331),
            .I(N__20317));
    LocalMux I__4818 (
            .O(N__20328),
            .I(N__20312));
    Span4Mux_h I__4817 (
            .O(N__20325),
            .I(N__20312));
    Span4Mux_v I__4816 (
            .O(N__20320),
            .I(N__20309));
    LocalMux I__4815 (
            .O(N__20317),
            .I(N__20303));
    Span4Mux_v I__4814 (
            .O(N__20312),
            .I(N__20303));
    Span4Mux_v I__4813 (
            .O(N__20309),
            .I(N__20300));
    InMux I__4812 (
            .O(N__20308),
            .I(N__20297));
    Span4Mux_v I__4811 (
            .O(N__20303),
            .I(N__20294));
    Span4Mux_v I__4810 (
            .O(N__20300),
            .I(N__20291));
    LocalMux I__4809 (
            .O(N__20297),
            .I(\Lab_UT.scctrl.next_state_0_2 ));
    Odrv4 I__4808 (
            .O(N__20294),
            .I(\Lab_UT.scctrl.next_state_0_2 ));
    Odrv4 I__4807 (
            .O(N__20291),
            .I(\Lab_UT.scctrl.next_state_0_2 ));
    InMux I__4806 (
            .O(N__20284),
            .I(N__20279));
    InMux I__4805 (
            .O(N__20283),
            .I(N__20276));
    CascadeMux I__4804 (
            .O(N__20282),
            .I(N__20273));
    LocalMux I__4803 (
            .O(N__20279),
            .I(N__20264));
    LocalMux I__4802 (
            .O(N__20276),
            .I(N__20261));
    InMux I__4801 (
            .O(N__20273),
            .I(N__20258));
    CascadeMux I__4800 (
            .O(N__20272),
            .I(N__20253));
    InMux I__4799 (
            .O(N__20271),
            .I(N__20250));
    InMux I__4798 (
            .O(N__20270),
            .I(N__20247));
    InMux I__4797 (
            .O(N__20269),
            .I(N__20244));
    InMux I__4796 (
            .O(N__20268),
            .I(N__20240));
    InMux I__4795 (
            .O(N__20267),
            .I(N__20237));
    Span4Mux_v I__4794 (
            .O(N__20264),
            .I(N__20230));
    Span4Mux_h I__4793 (
            .O(N__20261),
            .I(N__20230));
    LocalMux I__4792 (
            .O(N__20258),
            .I(N__20230));
    CascadeMux I__4791 (
            .O(N__20257),
            .I(N__20226));
    InMux I__4790 (
            .O(N__20256),
            .I(N__20223));
    InMux I__4789 (
            .O(N__20253),
            .I(N__20219));
    LocalMux I__4788 (
            .O(N__20250),
            .I(N__20216));
    LocalMux I__4787 (
            .O(N__20247),
            .I(N__20213));
    LocalMux I__4786 (
            .O(N__20244),
            .I(N__20210));
    InMux I__4785 (
            .O(N__20243),
            .I(N__20206));
    LocalMux I__4784 (
            .O(N__20240),
            .I(N__20201));
    LocalMux I__4783 (
            .O(N__20237),
            .I(N__20201));
    Span4Mux_v I__4782 (
            .O(N__20230),
            .I(N__20198));
    InMux I__4781 (
            .O(N__20229),
            .I(N__20195));
    InMux I__4780 (
            .O(N__20226),
            .I(N__20192));
    LocalMux I__4779 (
            .O(N__20223),
            .I(N__20189));
    CascadeMux I__4778 (
            .O(N__20222),
            .I(N__20185));
    LocalMux I__4777 (
            .O(N__20219),
            .I(N__20179));
    Span4Mux_v I__4776 (
            .O(N__20216),
            .I(N__20179));
    Span4Mux_v I__4775 (
            .O(N__20213),
            .I(N__20174));
    Span4Mux_s1_h I__4774 (
            .O(N__20210),
            .I(N__20174));
    InMux I__4773 (
            .O(N__20209),
            .I(N__20171));
    LocalMux I__4772 (
            .O(N__20206),
            .I(N__20168));
    Span4Mux_v I__4771 (
            .O(N__20201),
            .I(N__20165));
    Span4Mux_h I__4770 (
            .O(N__20198),
            .I(N__20156));
    LocalMux I__4769 (
            .O(N__20195),
            .I(N__20156));
    LocalMux I__4768 (
            .O(N__20192),
            .I(N__20156));
    Span4Mux_s3_v I__4767 (
            .O(N__20189),
            .I(N__20152));
    InMux I__4766 (
            .O(N__20188),
            .I(N__20147));
    InMux I__4765 (
            .O(N__20185),
            .I(N__20147));
    InMux I__4764 (
            .O(N__20184),
            .I(N__20144));
    Span4Mux_h I__4763 (
            .O(N__20179),
            .I(N__20137));
    Span4Mux_h I__4762 (
            .O(N__20174),
            .I(N__20137));
    LocalMux I__4761 (
            .O(N__20171),
            .I(N__20137));
    Span4Mux_h I__4760 (
            .O(N__20168),
            .I(N__20132));
    Span4Mux_v I__4759 (
            .O(N__20165),
            .I(N__20132));
    InMux I__4758 (
            .O(N__20164),
            .I(N__20127));
    InMux I__4757 (
            .O(N__20163),
            .I(N__20127));
    Span4Mux_h I__4756 (
            .O(N__20156),
            .I(N__20124));
    InMux I__4755 (
            .O(N__20155),
            .I(N__20121));
    Sp12to4 I__4754 (
            .O(N__20152),
            .I(N__20116));
    LocalMux I__4753 (
            .O(N__20147),
            .I(N__20116));
    LocalMux I__4752 (
            .O(N__20144),
            .I(N__20111));
    Span4Mux_v I__4751 (
            .O(N__20137),
            .I(N__20111));
    Odrv4 I__4750 (
            .O(N__20132),
            .I(rst_i_3));
    LocalMux I__4749 (
            .O(N__20127),
            .I(rst_i_3));
    Odrv4 I__4748 (
            .O(N__20124),
            .I(rst_i_3));
    LocalMux I__4747 (
            .O(N__20121),
            .I(rst_i_3));
    Odrv12 I__4746 (
            .O(N__20116),
            .I(rst_i_3));
    Odrv4 I__4745 (
            .O(N__20111),
            .I(rst_i_3));
    InMux I__4744 (
            .O(N__20098),
            .I(N__20085));
    CascadeMux I__4743 (
            .O(N__20097),
            .I(N__20072));
    InMux I__4742 (
            .O(N__20096),
            .I(N__20066));
    InMux I__4741 (
            .O(N__20095),
            .I(N__20063));
    CascadeMux I__4740 (
            .O(N__20094),
            .I(N__20056));
    CascadeMux I__4739 (
            .O(N__20093),
            .I(N__20053));
    InMux I__4738 (
            .O(N__20092),
            .I(N__20041));
    InMux I__4737 (
            .O(N__20091),
            .I(N__20041));
    InMux I__4736 (
            .O(N__20090),
            .I(N__20041));
    InMux I__4735 (
            .O(N__20089),
            .I(N__20041));
    InMux I__4734 (
            .O(N__20088),
            .I(N__20038));
    LocalMux I__4733 (
            .O(N__20085),
            .I(N__20035));
    InMux I__4732 (
            .O(N__20084),
            .I(N__20028));
    InMux I__4731 (
            .O(N__20083),
            .I(N__20028));
    InMux I__4730 (
            .O(N__20082),
            .I(N__20028));
    InMux I__4729 (
            .O(N__20081),
            .I(N__20021));
    InMux I__4728 (
            .O(N__20080),
            .I(N__20021));
    InMux I__4727 (
            .O(N__20079),
            .I(N__20021));
    InMux I__4726 (
            .O(N__20078),
            .I(N__20015));
    InMux I__4725 (
            .O(N__20077),
            .I(N__20012));
    InMux I__4724 (
            .O(N__20076),
            .I(N__20009));
    InMux I__4723 (
            .O(N__20075),
            .I(N__20002));
    InMux I__4722 (
            .O(N__20072),
            .I(N__20002));
    InMux I__4721 (
            .O(N__20071),
            .I(N__20002));
    InMux I__4720 (
            .O(N__20070),
            .I(N__19999));
    CascadeMux I__4719 (
            .O(N__20069),
            .I(N__19993));
    LocalMux I__4718 (
            .O(N__20066),
            .I(N__19987));
    LocalMux I__4717 (
            .O(N__20063),
            .I(N__19987));
    InMux I__4716 (
            .O(N__20062),
            .I(N__19984));
    InMux I__4715 (
            .O(N__20061),
            .I(N__19981));
    InMux I__4714 (
            .O(N__20060),
            .I(N__19978));
    InMux I__4713 (
            .O(N__20059),
            .I(N__19973));
    InMux I__4712 (
            .O(N__20056),
            .I(N__19973));
    InMux I__4711 (
            .O(N__20053),
            .I(N__19958));
    InMux I__4710 (
            .O(N__20052),
            .I(N__19955));
    InMux I__4709 (
            .O(N__20051),
            .I(N__19952));
    InMux I__4708 (
            .O(N__20050),
            .I(N__19949));
    LocalMux I__4707 (
            .O(N__20041),
            .I(N__19944));
    LocalMux I__4706 (
            .O(N__20038),
            .I(N__19944));
    Span4Mux_v I__4705 (
            .O(N__20035),
            .I(N__19941));
    LocalMux I__4704 (
            .O(N__20028),
            .I(N__19936));
    LocalMux I__4703 (
            .O(N__20021),
            .I(N__19936));
    InMux I__4702 (
            .O(N__20020),
            .I(N__19931));
    InMux I__4701 (
            .O(N__20019),
            .I(N__19931));
    InMux I__4700 (
            .O(N__20018),
            .I(N__19928));
    LocalMux I__4699 (
            .O(N__20015),
            .I(N__19923));
    LocalMux I__4698 (
            .O(N__20012),
            .I(N__19923));
    LocalMux I__4697 (
            .O(N__20009),
            .I(N__19918));
    LocalMux I__4696 (
            .O(N__20002),
            .I(N__19918));
    LocalMux I__4695 (
            .O(N__19999),
            .I(N__19912));
    InMux I__4694 (
            .O(N__19998),
            .I(N__19909));
    InMux I__4693 (
            .O(N__19997),
            .I(N__19904));
    InMux I__4692 (
            .O(N__19996),
            .I(N__19904));
    InMux I__4691 (
            .O(N__19993),
            .I(N__19899));
    InMux I__4690 (
            .O(N__19992),
            .I(N__19899));
    Span4Mux_v I__4689 (
            .O(N__19987),
            .I(N__19894));
    LocalMux I__4688 (
            .O(N__19984),
            .I(N__19894));
    LocalMux I__4687 (
            .O(N__19981),
            .I(N__19889));
    LocalMux I__4686 (
            .O(N__19978),
            .I(N__19889));
    LocalMux I__4685 (
            .O(N__19973),
            .I(N__19886));
    InMux I__4684 (
            .O(N__19972),
            .I(N__19881));
    InMux I__4683 (
            .O(N__19971),
            .I(N__19881));
    InMux I__4682 (
            .O(N__19970),
            .I(N__19872));
    InMux I__4681 (
            .O(N__19969),
            .I(N__19869));
    InMux I__4680 (
            .O(N__19968),
            .I(N__19866));
    InMux I__4679 (
            .O(N__19967),
            .I(N__19857));
    InMux I__4678 (
            .O(N__19966),
            .I(N__19857));
    InMux I__4677 (
            .O(N__19965),
            .I(N__19857));
    InMux I__4676 (
            .O(N__19964),
            .I(N__19857));
    InMux I__4675 (
            .O(N__19963),
            .I(N__19850));
    InMux I__4674 (
            .O(N__19962),
            .I(N__19850));
    InMux I__4673 (
            .O(N__19961),
            .I(N__19850));
    LocalMux I__4672 (
            .O(N__19958),
            .I(N__19847));
    LocalMux I__4671 (
            .O(N__19955),
            .I(N__19836));
    LocalMux I__4670 (
            .O(N__19952),
            .I(N__19836));
    LocalMux I__4669 (
            .O(N__19949),
            .I(N__19836));
    Span4Mux_v I__4668 (
            .O(N__19944),
            .I(N__19836));
    Span4Mux_h I__4667 (
            .O(N__19941),
            .I(N__19836));
    Span4Mux_h I__4666 (
            .O(N__19936),
            .I(N__19831));
    LocalMux I__4665 (
            .O(N__19931),
            .I(N__19828));
    LocalMux I__4664 (
            .O(N__19928),
            .I(N__19821));
    Span4Mux_v I__4663 (
            .O(N__19923),
            .I(N__19821));
    Span4Mux_v I__4662 (
            .O(N__19918),
            .I(N__19821));
    InMux I__4661 (
            .O(N__19917),
            .I(N__19814));
    InMux I__4660 (
            .O(N__19916),
            .I(N__19814));
    InMux I__4659 (
            .O(N__19915),
            .I(N__19814));
    Span4Mux_v I__4658 (
            .O(N__19912),
            .I(N__19807));
    LocalMux I__4657 (
            .O(N__19909),
            .I(N__19807));
    LocalMux I__4656 (
            .O(N__19904),
            .I(N__19807));
    LocalMux I__4655 (
            .O(N__19899),
            .I(N__19804));
    Span4Mux_h I__4654 (
            .O(N__19894),
            .I(N__19801));
    Span4Mux_h I__4653 (
            .O(N__19889),
            .I(N__19796));
    Span4Mux_v I__4652 (
            .O(N__19886),
            .I(N__19796));
    LocalMux I__4651 (
            .O(N__19881),
            .I(N__19793));
    InMux I__4650 (
            .O(N__19880),
            .I(N__19788));
    InMux I__4649 (
            .O(N__19879),
            .I(N__19788));
    InMux I__4648 (
            .O(N__19878),
            .I(N__19781));
    InMux I__4647 (
            .O(N__19877),
            .I(N__19781));
    InMux I__4646 (
            .O(N__19876),
            .I(N__19781));
    InMux I__4645 (
            .O(N__19875),
            .I(N__19778));
    LocalMux I__4644 (
            .O(N__19872),
            .I(N__19775));
    LocalMux I__4643 (
            .O(N__19869),
            .I(N__19762));
    LocalMux I__4642 (
            .O(N__19866),
            .I(N__19762));
    LocalMux I__4641 (
            .O(N__19857),
            .I(N__19762));
    LocalMux I__4640 (
            .O(N__19850),
            .I(N__19762));
    Span4Mux_v I__4639 (
            .O(N__19847),
            .I(N__19762));
    Span4Mux_v I__4638 (
            .O(N__19836),
            .I(N__19762));
    InMux I__4637 (
            .O(N__19835),
            .I(N__19757));
    InMux I__4636 (
            .O(N__19834),
            .I(N__19757));
    Span4Mux_v I__4635 (
            .O(N__19831),
            .I(N__19752));
    Span4Mux_s2_h I__4634 (
            .O(N__19828),
            .I(N__19752));
    Span4Mux_v I__4633 (
            .O(N__19821),
            .I(N__19743));
    LocalMux I__4632 (
            .O(N__19814),
            .I(N__19743));
    Span4Mux_v I__4631 (
            .O(N__19807),
            .I(N__19743));
    Span4Mux_v I__4630 (
            .O(N__19804),
            .I(N__19743));
    Span4Mux_v I__4629 (
            .O(N__19801),
            .I(N__19736));
    Span4Mux_v I__4628 (
            .O(N__19796),
            .I(N__19736));
    Span4Mux_s2_h I__4627 (
            .O(N__19793),
            .I(N__19736));
    LocalMux I__4626 (
            .O(N__19788),
            .I(Lab_UT_scctrl_N_221_0));
    LocalMux I__4625 (
            .O(N__19781),
            .I(Lab_UT_scctrl_N_221_0));
    LocalMux I__4624 (
            .O(N__19778),
            .I(Lab_UT_scctrl_N_221_0));
    Odrv12 I__4623 (
            .O(N__19775),
            .I(Lab_UT_scctrl_N_221_0));
    Odrv4 I__4622 (
            .O(N__19762),
            .I(Lab_UT_scctrl_N_221_0));
    LocalMux I__4621 (
            .O(N__19757),
            .I(Lab_UT_scctrl_N_221_0));
    Odrv4 I__4620 (
            .O(N__19752),
            .I(Lab_UT_scctrl_N_221_0));
    Odrv4 I__4619 (
            .O(N__19743),
            .I(Lab_UT_scctrl_N_221_0));
    Odrv4 I__4618 (
            .O(N__19736),
            .I(Lab_UT_scctrl_N_221_0));
    InMux I__4617 (
            .O(N__19717),
            .I(N__19711));
    InMux I__4616 (
            .O(N__19716),
            .I(N__19711));
    LocalMux I__4615 (
            .O(N__19711),
            .I(N__19708));
    Odrv12 I__4614 (
            .O(N__19708),
            .I(\Lab_UT.scctrl.G_21_i_0 ));
    InMux I__4613 (
            .O(N__19705),
            .I(N__19700));
    CascadeMux I__4612 (
            .O(N__19704),
            .I(N__19692));
    InMux I__4611 (
            .O(N__19703),
            .I(N__19688));
    LocalMux I__4610 (
            .O(N__19700),
            .I(N__19685));
    InMux I__4609 (
            .O(N__19699),
            .I(N__19680));
    InMux I__4608 (
            .O(N__19698),
            .I(N__19680));
    InMux I__4607 (
            .O(N__19697),
            .I(N__19675));
    InMux I__4606 (
            .O(N__19696),
            .I(N__19670));
    InMux I__4605 (
            .O(N__19695),
            .I(N__19670));
    InMux I__4604 (
            .O(N__19692),
            .I(N__19667));
    CascadeMux I__4603 (
            .O(N__19691),
            .I(N__19663));
    LocalMux I__4602 (
            .O(N__19688),
            .I(N__19659));
    Span4Mux_v I__4601 (
            .O(N__19685),
            .I(N__19655));
    LocalMux I__4600 (
            .O(N__19680),
            .I(N__19651));
    InMux I__4599 (
            .O(N__19679),
            .I(N__19646));
    InMux I__4598 (
            .O(N__19678),
            .I(N__19646));
    LocalMux I__4597 (
            .O(N__19675),
            .I(N__19643));
    LocalMux I__4596 (
            .O(N__19670),
            .I(N__19640));
    LocalMux I__4595 (
            .O(N__19667),
            .I(N__19637));
    InMux I__4594 (
            .O(N__19666),
            .I(N__19632));
    InMux I__4593 (
            .O(N__19663),
            .I(N__19632));
    InMux I__4592 (
            .O(N__19662),
            .I(N__19629));
    Span4Mux_h I__4591 (
            .O(N__19659),
            .I(N__19625));
    InMux I__4590 (
            .O(N__19658),
            .I(N__19622));
    IoSpan4Mux I__4589 (
            .O(N__19655),
            .I(N__19618));
    InMux I__4588 (
            .O(N__19654),
            .I(N__19615));
    Span4Mux_s3_v I__4587 (
            .O(N__19651),
            .I(N__19612));
    LocalMux I__4586 (
            .O(N__19646),
            .I(N__19605));
    Span4Mux_h I__4585 (
            .O(N__19643),
            .I(N__19605));
    Span4Mux_v I__4584 (
            .O(N__19640),
            .I(N__19605));
    Span4Mux_s2_v I__4583 (
            .O(N__19637),
            .I(N__19598));
    LocalMux I__4582 (
            .O(N__19632),
            .I(N__19598));
    LocalMux I__4581 (
            .O(N__19629),
            .I(N__19598));
    InMux I__4580 (
            .O(N__19628),
            .I(N__19595));
    Span4Mux_v I__4579 (
            .O(N__19625),
            .I(N__19592));
    LocalMux I__4578 (
            .O(N__19622),
            .I(N__19589));
    InMux I__4577 (
            .O(N__19621),
            .I(N__19586));
    Span4Mux_s1_h I__4576 (
            .O(N__19618),
            .I(N__19579));
    LocalMux I__4575 (
            .O(N__19615),
            .I(N__19579));
    Span4Mux_h I__4574 (
            .O(N__19612),
            .I(N__19579));
    Span4Mux_v I__4573 (
            .O(N__19605),
            .I(N__19574));
    Span4Mux_v I__4572 (
            .O(N__19598),
            .I(N__19574));
    LocalMux I__4571 (
            .O(N__19595),
            .I(\Lab_UT.state_i_3_2 ));
    Odrv4 I__4570 (
            .O(N__19592),
            .I(\Lab_UT.state_i_3_2 ));
    Odrv4 I__4569 (
            .O(N__19589),
            .I(\Lab_UT.state_i_3_2 ));
    LocalMux I__4568 (
            .O(N__19586),
            .I(\Lab_UT.state_i_3_2 ));
    Odrv4 I__4567 (
            .O(N__19579),
            .I(\Lab_UT.state_i_3_2 ));
    Odrv4 I__4566 (
            .O(N__19574),
            .I(\Lab_UT.state_i_3_2 ));
    CascadeMux I__4565 (
            .O(N__19561),
            .I(N__19557));
    InMux I__4564 (
            .O(N__19560),
            .I(N__19547));
    InMux I__4563 (
            .O(N__19557),
            .I(N__19544));
    InMux I__4562 (
            .O(N__19556),
            .I(N__19539));
    InMux I__4561 (
            .O(N__19555),
            .I(N__19539));
    CascadeMux I__4560 (
            .O(N__19554),
            .I(N__19534));
    CascadeMux I__4559 (
            .O(N__19553),
            .I(N__19531));
    InMux I__4558 (
            .O(N__19552),
            .I(N__19525));
    InMux I__4557 (
            .O(N__19551),
            .I(N__19525));
    CascadeMux I__4556 (
            .O(N__19550),
            .I(N__19522));
    LocalMux I__4555 (
            .O(N__19547),
            .I(N__19518));
    LocalMux I__4554 (
            .O(N__19544),
            .I(N__19515));
    LocalMux I__4553 (
            .O(N__19539),
            .I(N__19512));
    InMux I__4552 (
            .O(N__19538),
            .I(N__19509));
    InMux I__4551 (
            .O(N__19537),
            .I(N__19506));
    InMux I__4550 (
            .O(N__19534),
            .I(N__19503));
    InMux I__4549 (
            .O(N__19531),
            .I(N__19500));
    InMux I__4548 (
            .O(N__19530),
            .I(N__19497));
    LocalMux I__4547 (
            .O(N__19525),
            .I(N__19494));
    InMux I__4546 (
            .O(N__19522),
            .I(N__19491));
    InMux I__4545 (
            .O(N__19521),
            .I(N__19488));
    Span4Mux_v I__4544 (
            .O(N__19518),
            .I(N__19474));
    Span4Mux_h I__4543 (
            .O(N__19515),
            .I(N__19474));
    Span4Mux_v I__4542 (
            .O(N__19512),
            .I(N__19474));
    LocalMux I__4541 (
            .O(N__19509),
            .I(N__19474));
    LocalMux I__4540 (
            .O(N__19506),
            .I(N__19474));
    LocalMux I__4539 (
            .O(N__19503),
            .I(N__19471));
    LocalMux I__4538 (
            .O(N__19500),
            .I(N__19468));
    LocalMux I__4537 (
            .O(N__19497),
            .I(N__19463));
    Span4Mux_h I__4536 (
            .O(N__19494),
            .I(N__19463));
    LocalMux I__4535 (
            .O(N__19491),
            .I(N__19460));
    LocalMux I__4534 (
            .O(N__19488),
            .I(N__19457));
    InMux I__4533 (
            .O(N__19487),
            .I(N__19450));
    InMux I__4532 (
            .O(N__19486),
            .I(N__19450));
    InMux I__4531 (
            .O(N__19485),
            .I(N__19450));
    Span4Mux_h I__4530 (
            .O(N__19474),
            .I(N__19447));
    Span4Mux_v I__4529 (
            .O(N__19471),
            .I(N__19440));
    Span4Mux_h I__4528 (
            .O(N__19468),
            .I(N__19440));
    Span4Mux_v I__4527 (
            .O(N__19463),
            .I(N__19440));
    Odrv4 I__4526 (
            .O(N__19460),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__4525 (
            .O(N__19457),
            .I(\Lab_UT.state_2 ));
    LocalMux I__4524 (
            .O(N__19450),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__4523 (
            .O(N__19447),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__4522 (
            .O(N__19440),
            .I(\Lab_UT.state_2 ));
    InMux I__4521 (
            .O(N__19429),
            .I(N__19426));
    LocalMux I__4520 (
            .O(N__19426),
            .I(N__19422));
    InMux I__4519 (
            .O(N__19425),
            .I(N__19419));
    Span4Mux_s2_h I__4518 (
            .O(N__19422),
            .I(N__19416));
    LocalMux I__4517 (
            .O(N__19419),
            .I(N__19413));
    Odrv4 I__4516 (
            .O(N__19416),
            .I(\Lab_UT.scctrl.N_11_1 ));
    Odrv4 I__4515 (
            .O(N__19413),
            .I(\Lab_UT.scctrl.N_11_1 ));
    InMux I__4514 (
            .O(N__19408),
            .I(N__19405));
    LocalMux I__4513 (
            .O(N__19405),
            .I(N__19402));
    Span4Mux_s3_h I__4512 (
            .O(N__19402),
            .I(N__19399));
    Odrv4 I__4511 (
            .O(N__19399),
            .I(\Lab_UT.scctrl.N_12_2 ));
    CascadeMux I__4510 (
            .O(N__19396),
            .I(\Lab_UT.scctrl.G_24_i_a4_1_cascade_ ));
    CascadeMux I__4509 (
            .O(N__19393),
            .I(N__19390));
    InMux I__4508 (
            .O(N__19390),
            .I(N__19387));
    LocalMux I__4507 (
            .O(N__19387),
            .I(N__19384));
    Odrv4 I__4506 (
            .O(N__19384),
            .I(\Lab_UT.scctrl.G_21_i_a7_0_1 ));
    InMux I__4505 (
            .O(N__19381),
            .I(N__19372));
    InMux I__4504 (
            .O(N__19380),
            .I(N__19372));
    InMux I__4503 (
            .O(N__19379),
            .I(N__19372));
    LocalMux I__4502 (
            .O(N__19372),
            .I(N__19368));
    InMux I__4501 (
            .O(N__19371),
            .I(N__19365));
    Odrv4 I__4500 (
            .O(N__19368),
            .I(\Lab_UT.scctrl.N_9_2 ));
    LocalMux I__4499 (
            .O(N__19365),
            .I(\Lab_UT.scctrl.N_9_2 ));
    CascadeMux I__4498 (
            .O(N__19360),
            .I(N__19356));
    CascadeMux I__4497 (
            .O(N__19359),
            .I(N__19353));
    InMux I__4496 (
            .O(N__19356),
            .I(N__19348));
    InMux I__4495 (
            .O(N__19353),
            .I(N__19348));
    LocalMux I__4494 (
            .O(N__19348),
            .I(\Lab_UT.scctrl.G_21_i_2 ));
    InMux I__4493 (
            .O(N__19345),
            .I(N__19335));
    InMux I__4492 (
            .O(N__19344),
            .I(N__19335));
    InMux I__4491 (
            .O(N__19343),
            .I(N__19335));
    InMux I__4490 (
            .O(N__19342),
            .I(N__19332));
    LocalMux I__4489 (
            .O(N__19335),
            .I(\Lab_UT.scctrl.N_8_2 ));
    LocalMux I__4488 (
            .O(N__19332),
            .I(\Lab_UT.scctrl.N_8_2 ));
    CascadeMux I__4487 (
            .O(N__19327),
            .I(N__19324));
    InMux I__4486 (
            .O(N__19324),
            .I(N__19320));
    CascadeMux I__4485 (
            .O(N__19323),
            .I(N__19316));
    LocalMux I__4484 (
            .O(N__19320),
            .I(N__19311));
    InMux I__4483 (
            .O(N__19319),
            .I(N__19306));
    InMux I__4482 (
            .O(N__19316),
            .I(N__19303));
    InMux I__4481 (
            .O(N__19315),
            .I(N__19300));
    InMux I__4480 (
            .O(N__19314),
            .I(N__19297));
    Span4Mux_s2_h I__4479 (
            .O(N__19311),
            .I(N__19294));
    InMux I__4478 (
            .O(N__19310),
            .I(N__19289));
    InMux I__4477 (
            .O(N__19309),
            .I(N__19286));
    LocalMux I__4476 (
            .O(N__19306),
            .I(N__19281));
    LocalMux I__4475 (
            .O(N__19303),
            .I(N__19281));
    LocalMux I__4474 (
            .O(N__19300),
            .I(N__19278));
    LocalMux I__4473 (
            .O(N__19297),
            .I(N__19275));
    Span4Mux_v I__4472 (
            .O(N__19294),
            .I(N__19272));
    InMux I__4471 (
            .O(N__19293),
            .I(N__19269));
    InMux I__4470 (
            .O(N__19292),
            .I(N__19266));
    LocalMux I__4469 (
            .O(N__19289),
            .I(N__19263));
    LocalMux I__4468 (
            .O(N__19286),
            .I(N__19254));
    Span4Mux_s3_h I__4467 (
            .O(N__19281),
            .I(N__19254));
    Span4Mux_v I__4466 (
            .O(N__19278),
            .I(N__19254));
    Span4Mux_v I__4465 (
            .O(N__19275),
            .I(N__19254));
    Odrv4 I__4464 (
            .O(N__19272),
            .I(\Lab_UT.state_i_3_0_rep1 ));
    LocalMux I__4463 (
            .O(N__19269),
            .I(\Lab_UT.state_i_3_0_rep1 ));
    LocalMux I__4462 (
            .O(N__19266),
            .I(\Lab_UT.state_i_3_0_rep1 ));
    Odrv4 I__4461 (
            .O(N__19263),
            .I(\Lab_UT.state_i_3_0_rep1 ));
    Odrv4 I__4460 (
            .O(N__19254),
            .I(\Lab_UT.state_i_3_0_rep1 ));
    InMux I__4459 (
            .O(N__19243),
            .I(N__19240));
    LocalMux I__4458 (
            .O(N__19240),
            .I(N__19234));
    InMux I__4457 (
            .O(N__19239),
            .I(N__19231));
    InMux I__4456 (
            .O(N__19238),
            .I(N__19228));
    InMux I__4455 (
            .O(N__19237),
            .I(N__19225));
    Span4Mux_v I__4454 (
            .O(N__19234),
            .I(N__19220));
    LocalMux I__4453 (
            .O(N__19231),
            .I(N__19220));
    LocalMux I__4452 (
            .O(N__19228),
            .I(N__19216));
    LocalMux I__4451 (
            .O(N__19225),
            .I(N__19213));
    Span4Mux_h I__4450 (
            .O(N__19220),
            .I(N__19207));
    InMux I__4449 (
            .O(N__19219),
            .I(N__19204));
    Span12Mux_s4_h I__4448 (
            .O(N__19216),
            .I(N__19199));
    Span12Mux_s5_v I__4447 (
            .O(N__19213),
            .I(N__19199));
    InMux I__4446 (
            .O(N__19212),
            .I(N__19194));
    InMux I__4445 (
            .O(N__19211),
            .I(N__19194));
    InMux I__4444 (
            .O(N__19210),
            .I(N__19191));
    Odrv4 I__4443 (
            .O(N__19207),
            .I(\Lab_UT.state_i_3_2_rep1 ));
    LocalMux I__4442 (
            .O(N__19204),
            .I(\Lab_UT.state_i_3_2_rep1 ));
    Odrv12 I__4441 (
            .O(N__19199),
            .I(\Lab_UT.state_i_3_2_rep1 ));
    LocalMux I__4440 (
            .O(N__19194),
            .I(\Lab_UT.state_i_3_2_rep1 ));
    LocalMux I__4439 (
            .O(N__19191),
            .I(\Lab_UT.state_i_3_2_rep1 ));
    InMux I__4438 (
            .O(N__19180),
            .I(N__19177));
    LocalMux I__4437 (
            .O(N__19177),
            .I(N__19174));
    Odrv4 I__4436 (
            .O(N__19174),
            .I(\Lab_UT.scctrl.g0_1_4_1 ));
    CascadeMux I__4435 (
            .O(N__19171),
            .I(\Lab_UT.scctrl.g0_i_a7_0_1_cascade_ ));
    InMux I__4434 (
            .O(N__19168),
            .I(N__19158));
    CascadeMux I__4433 (
            .O(N__19167),
            .I(N__19152));
    InMux I__4432 (
            .O(N__19166),
            .I(N__19144));
    InMux I__4431 (
            .O(N__19165),
            .I(N__19139));
    InMux I__4430 (
            .O(N__19164),
            .I(N__19139));
    InMux I__4429 (
            .O(N__19163),
            .I(N__19134));
    InMux I__4428 (
            .O(N__19162),
            .I(N__19134));
    InMux I__4427 (
            .O(N__19161),
            .I(N__19131));
    LocalMux I__4426 (
            .O(N__19158),
            .I(N__19128));
    InMux I__4425 (
            .O(N__19157),
            .I(N__19125));
    InMux I__4424 (
            .O(N__19156),
            .I(N__19122));
    InMux I__4423 (
            .O(N__19155),
            .I(N__19119));
    InMux I__4422 (
            .O(N__19152),
            .I(N__19113));
    InMux I__4421 (
            .O(N__19151),
            .I(N__19113));
    InMux I__4420 (
            .O(N__19150),
            .I(N__19110));
    InMux I__4419 (
            .O(N__19149),
            .I(N__19102));
    InMux I__4418 (
            .O(N__19148),
            .I(N__19102));
    InMux I__4417 (
            .O(N__19147),
            .I(N__19098));
    LocalMux I__4416 (
            .O(N__19144),
            .I(N__19091));
    LocalMux I__4415 (
            .O(N__19139),
            .I(N__19091));
    LocalMux I__4414 (
            .O(N__19134),
            .I(N__19087));
    LocalMux I__4413 (
            .O(N__19131),
            .I(N__19084));
    Span4Mux_v I__4412 (
            .O(N__19128),
            .I(N__19079));
    LocalMux I__4411 (
            .O(N__19125),
            .I(N__19079));
    LocalMux I__4410 (
            .O(N__19122),
            .I(N__19076));
    LocalMux I__4409 (
            .O(N__19119),
            .I(N__19073));
    CascadeMux I__4408 (
            .O(N__19118),
            .I(N__19070));
    LocalMux I__4407 (
            .O(N__19113),
            .I(N__19066));
    LocalMux I__4406 (
            .O(N__19110),
            .I(N__19063));
    InMux I__4405 (
            .O(N__19109),
            .I(N__19058));
    InMux I__4404 (
            .O(N__19108),
            .I(N__19058));
    InMux I__4403 (
            .O(N__19107),
            .I(N__19055));
    LocalMux I__4402 (
            .O(N__19102),
            .I(N__19052));
    InMux I__4401 (
            .O(N__19101),
            .I(N__19049));
    LocalMux I__4400 (
            .O(N__19098),
            .I(N__19046));
    InMux I__4399 (
            .O(N__19097),
            .I(N__19041));
    InMux I__4398 (
            .O(N__19096),
            .I(N__19041));
    Span4Mux_h I__4397 (
            .O(N__19091),
            .I(N__19038));
    InMux I__4396 (
            .O(N__19090),
            .I(N__19035));
    Span4Mux_v I__4395 (
            .O(N__19087),
            .I(N__19032));
    Span4Mux_h I__4394 (
            .O(N__19084),
            .I(N__19027));
    Span4Mux_h I__4393 (
            .O(N__19079),
            .I(N__19027));
    Span4Mux_v I__4392 (
            .O(N__19076),
            .I(N__19022));
    Span4Mux_s1_h I__4391 (
            .O(N__19073),
            .I(N__19022));
    InMux I__4390 (
            .O(N__19070),
            .I(N__19017));
    InMux I__4389 (
            .O(N__19069),
            .I(N__19017));
    Span12Mux_s5_h I__4388 (
            .O(N__19066),
            .I(N__19010));
    Sp12to4 I__4387 (
            .O(N__19063),
            .I(N__19010));
    LocalMux I__4386 (
            .O(N__19058),
            .I(N__19010));
    LocalMux I__4385 (
            .O(N__19055),
            .I(N__19003));
    Span4Mux_h I__4384 (
            .O(N__19052),
            .I(N__19003));
    LocalMux I__4383 (
            .O(N__19049),
            .I(N__19003));
    Odrv4 I__4382 (
            .O(N__19046),
            .I(\Lab_UT.de_hex_0 ));
    LocalMux I__4381 (
            .O(N__19041),
            .I(\Lab_UT.de_hex_0 ));
    Odrv4 I__4380 (
            .O(N__19038),
            .I(\Lab_UT.de_hex_0 ));
    LocalMux I__4379 (
            .O(N__19035),
            .I(\Lab_UT.de_hex_0 ));
    Odrv4 I__4378 (
            .O(N__19032),
            .I(\Lab_UT.de_hex_0 ));
    Odrv4 I__4377 (
            .O(N__19027),
            .I(\Lab_UT.de_hex_0 ));
    Odrv4 I__4376 (
            .O(N__19022),
            .I(\Lab_UT.de_hex_0 ));
    LocalMux I__4375 (
            .O(N__19017),
            .I(\Lab_UT.de_hex_0 ));
    Odrv12 I__4374 (
            .O(N__19010),
            .I(\Lab_UT.de_hex_0 ));
    Odrv4 I__4373 (
            .O(N__19003),
            .I(\Lab_UT.de_hex_0 ));
    InMux I__4372 (
            .O(N__18982),
            .I(N__18979));
    LocalMux I__4371 (
            .O(N__18979),
            .I(N__18976));
    Odrv12 I__4370 (
            .O(N__18976),
            .I(\Lab_UT.scctrl.N_10_0 ));
    CascadeMux I__4369 (
            .O(N__18973),
            .I(\Lab_UT.scctrl.g0_7_a13_1_1_cascade_ ));
    CascadeMux I__4368 (
            .O(N__18970),
            .I(\Lab_UT.scctrl.N_7_cascade_ ));
    InMux I__4367 (
            .O(N__18967),
            .I(N__18964));
    LocalMux I__4366 (
            .O(N__18964),
            .I(N__18961));
    Span4Mux_h I__4365 (
            .O(N__18961),
            .I(N__18958));
    Odrv4 I__4364 (
            .O(N__18958),
            .I(\Lab_UT.scctrl.g0_6 ));
    InMux I__4363 (
            .O(N__18955),
            .I(N__18948));
    CascadeMux I__4362 (
            .O(N__18954),
            .I(N__18943));
    InMux I__4361 (
            .O(N__18953),
            .I(N__18940));
    InMux I__4360 (
            .O(N__18952),
            .I(N__18935));
    InMux I__4359 (
            .O(N__18951),
            .I(N__18932));
    LocalMux I__4358 (
            .O(N__18948),
            .I(N__18929));
    InMux I__4357 (
            .O(N__18947),
            .I(N__18926));
    InMux I__4356 (
            .O(N__18946),
            .I(N__18923));
    InMux I__4355 (
            .O(N__18943),
            .I(N__18919));
    LocalMux I__4354 (
            .O(N__18940),
            .I(N__18915));
    InMux I__4353 (
            .O(N__18939),
            .I(N__18910));
    InMux I__4352 (
            .O(N__18938),
            .I(N__18907));
    LocalMux I__4351 (
            .O(N__18935),
            .I(N__18904));
    LocalMux I__4350 (
            .O(N__18932),
            .I(N__18899));
    Span4Mux_s3_v I__4349 (
            .O(N__18929),
            .I(N__18899));
    LocalMux I__4348 (
            .O(N__18926),
            .I(N__18896));
    LocalMux I__4347 (
            .O(N__18923),
            .I(N__18893));
    InMux I__4346 (
            .O(N__18922),
            .I(N__18890));
    LocalMux I__4345 (
            .O(N__18919),
            .I(N__18887));
    InMux I__4344 (
            .O(N__18918),
            .I(N__18884));
    Span4Mux_s2_v I__4343 (
            .O(N__18915),
            .I(N__18881));
    InMux I__4342 (
            .O(N__18914),
            .I(N__18876));
    InMux I__4341 (
            .O(N__18913),
            .I(N__18876));
    LocalMux I__4340 (
            .O(N__18910),
            .I(N__18873));
    LocalMux I__4339 (
            .O(N__18907),
            .I(N__18870));
    Span4Mux_h I__4338 (
            .O(N__18904),
            .I(N__18864));
    Span4Mux_h I__4337 (
            .O(N__18899),
            .I(N__18864));
    Span4Mux_v I__4336 (
            .O(N__18896),
            .I(N__18859));
    Span4Mux_h I__4335 (
            .O(N__18893),
            .I(N__18859));
    LocalMux I__4334 (
            .O(N__18890),
            .I(N__18855));
    Span4Mux_v I__4333 (
            .O(N__18887),
            .I(N__18844));
    LocalMux I__4332 (
            .O(N__18884),
            .I(N__18844));
    Span4Mux_v I__4331 (
            .O(N__18881),
            .I(N__18844));
    LocalMux I__4330 (
            .O(N__18876),
            .I(N__18844));
    Span4Mux_v I__4329 (
            .O(N__18873),
            .I(N__18844));
    Span4Mux_s2_v I__4328 (
            .O(N__18870),
            .I(N__18841));
    InMux I__4327 (
            .O(N__18869),
            .I(N__18838));
    Span4Mux_v I__4326 (
            .O(N__18864),
            .I(N__18833));
    Span4Mux_h I__4325 (
            .O(N__18859),
            .I(N__18833));
    InMux I__4324 (
            .O(N__18858),
            .I(N__18830));
    Span4Mux_v I__4323 (
            .O(N__18855),
            .I(N__18823));
    Span4Mux_h I__4322 (
            .O(N__18844),
            .I(N__18823));
    Span4Mux_v I__4321 (
            .O(N__18841),
            .I(N__18823));
    LocalMux I__4320 (
            .O(N__18838),
            .I(rst));
    Odrv4 I__4319 (
            .O(N__18833),
            .I(rst));
    LocalMux I__4318 (
            .O(N__18830),
            .I(rst));
    Odrv4 I__4317 (
            .O(N__18823),
            .I(rst));
    InMux I__4316 (
            .O(N__18814),
            .I(N__18811));
    LocalMux I__4315 (
            .O(N__18811),
            .I(N__18808));
    Odrv12 I__4314 (
            .O(N__18808),
            .I(\Lab_UT.scctrl.g1_i_a7_2Z0Z_3 ));
    CascadeMux I__4313 (
            .O(N__18805),
            .I(\Lab_UT.scctrl.N_10_1_cascade_ ));
    InMux I__4312 (
            .O(N__18802),
            .I(N__18799));
    LocalMux I__4311 (
            .O(N__18799),
            .I(N__18796));
    Span4Mux_v I__4310 (
            .O(N__18796),
            .I(N__18793));
    Odrv4 I__4309 (
            .O(N__18793),
            .I(\Lab_UT.scctrl.g1_i_2 ));
    InMux I__4308 (
            .O(N__18790),
            .I(N__18787));
    LocalMux I__4307 (
            .O(N__18787),
            .I(\Lab_UT.scctrl.N_7_4 ));
    InMux I__4306 (
            .O(N__18784),
            .I(N__18777));
    InMux I__4305 (
            .O(N__18783),
            .I(N__18774));
    InMux I__4304 (
            .O(N__18782),
            .I(N__18766));
    InMux I__4303 (
            .O(N__18781),
            .I(N__18766));
    InMux I__4302 (
            .O(N__18780),
            .I(N__18760));
    LocalMux I__4301 (
            .O(N__18777),
            .I(N__18755));
    LocalMux I__4300 (
            .O(N__18774),
            .I(N__18755));
    InMux I__4299 (
            .O(N__18773),
            .I(N__18752));
    InMux I__4298 (
            .O(N__18772),
            .I(N__18745));
    InMux I__4297 (
            .O(N__18771),
            .I(N__18742));
    LocalMux I__4296 (
            .O(N__18766),
            .I(N__18739));
    InMux I__4295 (
            .O(N__18765),
            .I(N__18736));
    InMux I__4294 (
            .O(N__18764),
            .I(N__18731));
    InMux I__4293 (
            .O(N__18763),
            .I(N__18731));
    LocalMux I__4292 (
            .O(N__18760),
            .I(N__18725));
    Span4Mux_s3_h I__4291 (
            .O(N__18755),
            .I(N__18722));
    LocalMux I__4290 (
            .O(N__18752),
            .I(N__18716));
    InMux I__4289 (
            .O(N__18751),
            .I(N__18709));
    InMux I__4288 (
            .O(N__18750),
            .I(N__18709));
    InMux I__4287 (
            .O(N__18749),
            .I(N__18709));
    InMux I__4286 (
            .O(N__18748),
            .I(N__18706));
    LocalMux I__4285 (
            .O(N__18745),
            .I(N__18703));
    LocalMux I__4284 (
            .O(N__18742),
            .I(N__18698));
    Span4Mux_s3_v I__4283 (
            .O(N__18739),
            .I(N__18698));
    LocalMux I__4282 (
            .O(N__18736),
            .I(N__18695));
    LocalMux I__4281 (
            .O(N__18731),
            .I(N__18692));
    InMux I__4280 (
            .O(N__18730),
            .I(N__18689));
    InMux I__4279 (
            .O(N__18729),
            .I(N__18684));
    InMux I__4278 (
            .O(N__18728),
            .I(N__18684));
    Span4Mux_s3_h I__4277 (
            .O(N__18725),
            .I(N__18679));
    Span4Mux_v I__4276 (
            .O(N__18722),
            .I(N__18679));
    InMux I__4275 (
            .O(N__18721),
            .I(N__18672));
    InMux I__4274 (
            .O(N__18720),
            .I(N__18672));
    InMux I__4273 (
            .O(N__18719),
            .I(N__18672));
    Span4Mux_h I__4272 (
            .O(N__18716),
            .I(N__18667));
    LocalMux I__4271 (
            .O(N__18709),
            .I(N__18667));
    LocalMux I__4270 (
            .O(N__18706),
            .I(N__18658));
    Span4Mux_v I__4269 (
            .O(N__18703),
            .I(N__18658));
    Span4Mux_v I__4268 (
            .O(N__18698),
            .I(N__18658));
    Span4Mux_h I__4267 (
            .O(N__18695),
            .I(N__18658));
    Odrv12 I__4266 (
            .O(N__18692),
            .I(\Lab_UT.un1_de_hex ));
    LocalMux I__4265 (
            .O(N__18689),
            .I(\Lab_UT.un1_de_hex ));
    LocalMux I__4264 (
            .O(N__18684),
            .I(\Lab_UT.un1_de_hex ));
    Odrv4 I__4263 (
            .O(N__18679),
            .I(\Lab_UT.un1_de_hex ));
    LocalMux I__4262 (
            .O(N__18672),
            .I(\Lab_UT.un1_de_hex ));
    Odrv4 I__4261 (
            .O(N__18667),
            .I(\Lab_UT.un1_de_hex ));
    Odrv4 I__4260 (
            .O(N__18658),
            .I(\Lab_UT.un1_de_hex ));
    CascadeMux I__4259 (
            .O(N__18643),
            .I(N__18640));
    InMux I__4258 (
            .O(N__18640),
            .I(N__18637));
    LocalMux I__4257 (
            .O(N__18637),
            .I(N__18634));
    Span4Mux_s3_h I__4256 (
            .O(N__18634),
            .I(N__18631));
    Odrv4 I__4255 (
            .O(N__18631),
            .I(\Lab_UT.scctrl.G_21_i_a7_0 ));
    InMux I__4254 (
            .O(N__18628),
            .I(N__18617));
    CascadeMux I__4253 (
            .O(N__18627),
            .I(N__18613));
    InMux I__4252 (
            .O(N__18626),
            .I(N__18608));
    InMux I__4251 (
            .O(N__18625),
            .I(N__18605));
    InMux I__4250 (
            .O(N__18624),
            .I(N__18602));
    InMux I__4249 (
            .O(N__18623),
            .I(N__18592));
    InMux I__4248 (
            .O(N__18622),
            .I(N__18592));
    InMux I__4247 (
            .O(N__18621),
            .I(N__18592));
    InMux I__4246 (
            .O(N__18620),
            .I(N__18586));
    LocalMux I__4245 (
            .O(N__18617),
            .I(N__18583));
    InMux I__4244 (
            .O(N__18616),
            .I(N__18580));
    InMux I__4243 (
            .O(N__18613),
            .I(N__18573));
    InMux I__4242 (
            .O(N__18612),
            .I(N__18573));
    InMux I__4241 (
            .O(N__18611),
            .I(N__18573));
    LocalMux I__4240 (
            .O(N__18608),
            .I(N__18566));
    LocalMux I__4239 (
            .O(N__18605),
            .I(N__18566));
    LocalMux I__4238 (
            .O(N__18602),
            .I(N__18563));
    CascadeMux I__4237 (
            .O(N__18601),
            .I(N__18559));
    CascadeMux I__4236 (
            .O(N__18600),
            .I(N__18556));
    InMux I__4235 (
            .O(N__18599),
            .I(N__18553));
    LocalMux I__4234 (
            .O(N__18592),
            .I(N__18550));
    InMux I__4233 (
            .O(N__18591),
            .I(N__18547));
    CascadeMux I__4232 (
            .O(N__18590),
            .I(N__18544));
    CascadeMux I__4231 (
            .O(N__18589),
            .I(N__18540));
    LocalMux I__4230 (
            .O(N__18586),
            .I(N__18537));
    Span4Mux_v I__4229 (
            .O(N__18583),
            .I(N__18532));
    LocalMux I__4228 (
            .O(N__18580),
            .I(N__18532));
    LocalMux I__4227 (
            .O(N__18573),
            .I(N__18529));
    InMux I__4226 (
            .O(N__18572),
            .I(N__18524));
    InMux I__4225 (
            .O(N__18571),
            .I(N__18524));
    Span4Mux_v I__4224 (
            .O(N__18566),
            .I(N__18519));
    Span4Mux_v I__4223 (
            .O(N__18563),
            .I(N__18519));
    InMux I__4222 (
            .O(N__18562),
            .I(N__18512));
    InMux I__4221 (
            .O(N__18559),
            .I(N__18512));
    InMux I__4220 (
            .O(N__18556),
            .I(N__18512));
    LocalMux I__4219 (
            .O(N__18553),
            .I(N__18507));
    Span4Mux_v I__4218 (
            .O(N__18550),
            .I(N__18507));
    LocalMux I__4217 (
            .O(N__18547),
            .I(N__18504));
    InMux I__4216 (
            .O(N__18544),
            .I(N__18497));
    InMux I__4215 (
            .O(N__18543),
            .I(N__18497));
    InMux I__4214 (
            .O(N__18540),
            .I(N__18497));
    Span4Mux_h I__4213 (
            .O(N__18537),
            .I(N__18494));
    Span4Mux_h I__4212 (
            .O(N__18532),
            .I(N__18491));
    Odrv4 I__4211 (
            .O(N__18529),
            .I(\Lab_UT.un4_de_hex ));
    LocalMux I__4210 (
            .O(N__18524),
            .I(\Lab_UT.un4_de_hex ));
    Odrv4 I__4209 (
            .O(N__18519),
            .I(\Lab_UT.un4_de_hex ));
    LocalMux I__4208 (
            .O(N__18512),
            .I(\Lab_UT.un4_de_hex ));
    Odrv4 I__4207 (
            .O(N__18507),
            .I(\Lab_UT.un4_de_hex ));
    Odrv4 I__4206 (
            .O(N__18504),
            .I(\Lab_UT.un4_de_hex ));
    LocalMux I__4205 (
            .O(N__18497),
            .I(\Lab_UT.un4_de_hex ));
    Odrv4 I__4204 (
            .O(N__18494),
            .I(\Lab_UT.un4_de_hex ));
    Odrv4 I__4203 (
            .O(N__18491),
            .I(\Lab_UT.un4_de_hex ));
    CascadeMux I__4202 (
            .O(N__18472),
            .I(\Lab_UT.scctrl.g0_0_i_a8_0_1_cascade_ ));
    InMux I__4201 (
            .O(N__18469),
            .I(N__18466));
    LocalMux I__4200 (
            .O(N__18466),
            .I(N__18463));
    Span4Mux_v I__4199 (
            .O(N__18463),
            .I(N__18460));
    Span4Mux_h I__4198 (
            .O(N__18460),
            .I(N__18457));
    Odrv4 I__4197 (
            .O(N__18457),
            .I(\Lab_UT.scctrl.N_20 ));
    CascadeMux I__4196 (
            .O(N__18454),
            .I(\Lab_UT.scctrl.G_38_0_a3_0_4_cascade_ ));
    InMux I__4195 (
            .O(N__18451),
            .I(N__18447));
    CascadeMux I__4194 (
            .O(N__18450),
            .I(N__18444));
    LocalMux I__4193 (
            .O(N__18447),
            .I(N__18438));
    InMux I__4192 (
            .O(N__18444),
            .I(N__18435));
    CascadeMux I__4191 (
            .O(N__18443),
            .I(N__18432));
    InMux I__4190 (
            .O(N__18442),
            .I(N__18429));
    InMux I__4189 (
            .O(N__18441),
            .I(N__18426));
    Span4Mux_s1_h I__4188 (
            .O(N__18438),
            .I(N__18423));
    LocalMux I__4187 (
            .O(N__18435),
            .I(N__18419));
    InMux I__4186 (
            .O(N__18432),
            .I(N__18416));
    LocalMux I__4185 (
            .O(N__18429),
            .I(N__18413));
    LocalMux I__4184 (
            .O(N__18426),
            .I(N__18410));
    Span4Mux_v I__4183 (
            .O(N__18423),
            .I(N__18407));
    InMux I__4182 (
            .O(N__18422),
            .I(N__18404));
    Span4Mux_s3_v I__4181 (
            .O(N__18419),
            .I(N__18399));
    LocalMux I__4180 (
            .O(N__18416),
            .I(N__18399));
    Span12Mux_s9_v I__4179 (
            .O(N__18413),
            .I(N__18396));
    Span12Mux_s7_h I__4178 (
            .O(N__18410),
            .I(N__18393));
    Odrv4 I__4177 (
            .O(N__18407),
            .I(\Lab_UT.scctrl.next_stateZ0Z_0 ));
    LocalMux I__4176 (
            .O(N__18404),
            .I(\Lab_UT.scctrl.next_stateZ0Z_0 ));
    Odrv4 I__4175 (
            .O(N__18399),
            .I(\Lab_UT.scctrl.next_stateZ0Z_0 ));
    Odrv12 I__4174 (
            .O(N__18396),
            .I(\Lab_UT.scctrl.next_stateZ0Z_0 ));
    Odrv12 I__4173 (
            .O(N__18393),
            .I(\Lab_UT.scctrl.next_stateZ0Z_0 ));
    CascadeMux I__4172 (
            .O(N__18382),
            .I(\Lab_UT.scctrl.G_38_0_1_cascade_ ));
    InMux I__4171 (
            .O(N__18379),
            .I(N__18376));
    LocalMux I__4170 (
            .O(N__18376),
            .I(\Lab_UT.scctrl.N_7_0 ));
    InMux I__4169 (
            .O(N__18373),
            .I(N__18370));
    LocalMux I__4168 (
            .O(N__18370),
            .I(\Lab_UT.scctrl.g0_0_i_0 ));
    InMux I__4167 (
            .O(N__18367),
            .I(N__18364));
    LocalMux I__4166 (
            .O(N__18364),
            .I(N__18361));
    Odrv4 I__4165 (
            .O(N__18361),
            .I(\Lab_UT.scdp.a2b.g0_i_a9_1 ));
    CascadeMux I__4164 (
            .O(N__18358),
            .I(\Lab_UT.scdp.a2b.g0_iZ0Z_1_cascade_ ));
    InMux I__4163 (
            .O(N__18355),
            .I(N__18352));
    LocalMux I__4162 (
            .O(N__18352),
            .I(N__18349));
    Odrv12 I__4161 (
            .O(N__18349),
            .I(\Lab_UT.scdp.a2b.g0_iZ0Z_2 ));
    InMux I__4160 (
            .O(N__18346),
            .I(N__18343));
    LocalMux I__4159 (
            .O(N__18343),
            .I(N__18340));
    Odrv4 I__4158 (
            .O(N__18340),
            .I(\Lab_UT.scctrl.g1_i_a7_1 ));
    CascadeMux I__4157 (
            .O(N__18337),
            .I(N__18333));
    CascadeMux I__4156 (
            .O(N__18336),
            .I(N__18328));
    InMux I__4155 (
            .O(N__18333),
            .I(N__18322));
    CascadeMux I__4154 (
            .O(N__18332),
            .I(N__18319));
    CascadeMux I__4153 (
            .O(N__18331),
            .I(N__18316));
    InMux I__4152 (
            .O(N__18328),
            .I(N__18310));
    InMux I__4151 (
            .O(N__18327),
            .I(N__18310));
    InMux I__4150 (
            .O(N__18326),
            .I(N__18306));
    InMux I__4149 (
            .O(N__18325),
            .I(N__18303));
    LocalMux I__4148 (
            .O(N__18322),
            .I(N__18300));
    InMux I__4147 (
            .O(N__18319),
            .I(N__18293));
    InMux I__4146 (
            .O(N__18316),
            .I(N__18293));
    InMux I__4145 (
            .O(N__18315),
            .I(N__18293));
    LocalMux I__4144 (
            .O(N__18310),
            .I(N__18290));
    InMux I__4143 (
            .O(N__18309),
            .I(N__18287));
    LocalMux I__4142 (
            .O(N__18306),
            .I(N__18284));
    LocalMux I__4141 (
            .O(N__18303),
            .I(N__18281));
    Span4Mux_h I__4140 (
            .O(N__18300),
            .I(N__18276));
    LocalMux I__4139 (
            .O(N__18293),
            .I(N__18276));
    Span4Mux_h I__4138 (
            .O(N__18290),
            .I(N__18273));
    LocalMux I__4137 (
            .O(N__18287),
            .I(N__18270));
    Span4Mux_v I__4136 (
            .O(N__18284),
            .I(N__18263));
    Span4Mux_h I__4135 (
            .O(N__18281),
            .I(N__18263));
    Span4Mux_v I__4134 (
            .O(N__18276),
            .I(N__18263));
    Span4Mux_v I__4133 (
            .O(N__18273),
            .I(N__18260));
    Span4Mux_h I__4132 (
            .O(N__18270),
            .I(N__18257));
    Span4Mux_h I__4131 (
            .O(N__18263),
            .I(N__18254));
    Odrv4 I__4130 (
            .O(N__18260),
            .I(\Lab_UT.scctrl.next_state_0_3 ));
    Odrv4 I__4129 (
            .O(N__18257),
            .I(\Lab_UT.scctrl.next_state_0_3 ));
    Odrv4 I__4128 (
            .O(N__18254),
            .I(\Lab_UT.scctrl.next_state_0_3 ));
    InMux I__4127 (
            .O(N__18247),
            .I(N__18243));
    InMux I__4126 (
            .O(N__18246),
            .I(N__18240));
    LocalMux I__4125 (
            .O(N__18243),
            .I(N__18237));
    LocalMux I__4124 (
            .O(N__18240),
            .I(N__18231));
    Span4Mux_v I__4123 (
            .O(N__18237),
            .I(N__18231));
    InMux I__4122 (
            .O(N__18236),
            .I(N__18228));
    Odrv4 I__4121 (
            .O(N__18231),
            .I(\Lab_UT.scctrl.next_state_1_0_3 ));
    LocalMux I__4120 (
            .O(N__18228),
            .I(\Lab_UT.scctrl.next_state_1_0_3 ));
    CascadeMux I__4119 (
            .O(N__18223),
            .I(\Lab_UT.scctrl.next_state_i_3_cascade_ ));
    InMux I__4118 (
            .O(N__18220),
            .I(N__18217));
    LocalMux I__4117 (
            .O(N__18217),
            .I(N__18213));
    InMux I__4116 (
            .O(N__18216),
            .I(N__18210));
    Span4Mux_s3_v I__4115 (
            .O(N__18213),
            .I(N__18207));
    LocalMux I__4114 (
            .O(N__18210),
            .I(N__18204));
    Odrv4 I__4113 (
            .O(N__18207),
            .I(\Lab_UT.scctrl.next_state71 ));
    Odrv4 I__4112 (
            .O(N__18204),
            .I(\Lab_UT.scctrl.next_state71 ));
    InMux I__4111 (
            .O(N__18199),
            .I(N__18195));
    InMux I__4110 (
            .O(N__18198),
            .I(N__18192));
    LocalMux I__4109 (
            .O(N__18195),
            .I(N__18189));
    LocalMux I__4108 (
            .O(N__18192),
            .I(N__18186));
    Span4Mux_s3_v I__4107 (
            .O(N__18189),
            .I(N__18183));
    Span4Mux_h I__4106 (
            .O(N__18186),
            .I(N__18180));
    Odrv4 I__4105 (
            .O(N__18183),
            .I(\Lab_UT.scctrl.next_state72 ));
    Odrv4 I__4104 (
            .O(N__18180),
            .I(\Lab_UT.scctrl.next_state72 ));
    InMux I__4103 (
            .O(N__18175),
            .I(N__18172));
    LocalMux I__4102 (
            .O(N__18172),
            .I(N__18169));
    Odrv12 I__4101 (
            .O(N__18169),
            .I(\Lab_UT.scctrl.g4_1 ));
    InMux I__4100 (
            .O(N__18166),
            .I(N__18157));
    InMux I__4099 (
            .O(N__18165),
            .I(N__18157));
    InMux I__4098 (
            .O(N__18164),
            .I(N__18157));
    LocalMux I__4097 (
            .O(N__18157),
            .I(N__18152));
    InMux I__4096 (
            .O(N__18156),
            .I(N__18147));
    InMux I__4095 (
            .O(N__18155),
            .I(N__18147));
    Span4Mux_v I__4094 (
            .O(N__18152),
            .I(N__18142));
    LocalMux I__4093 (
            .O(N__18147),
            .I(N__18142));
    Span4Mux_v I__4092 (
            .O(N__18142),
            .I(N__18137));
    InMux I__4091 (
            .O(N__18141),
            .I(N__18134));
    InMux I__4090 (
            .O(N__18140),
            .I(N__18131));
    Span4Mux_h I__4089 (
            .O(N__18137),
            .I(N__18128));
    LocalMux I__4088 (
            .O(N__18134),
            .I(N__18125));
    LocalMux I__4087 (
            .O(N__18131),
            .I(\Lab_UT.sccEmsBitsSl ));
    Odrv4 I__4086 (
            .O(N__18128),
            .I(\Lab_UT.sccEmsBitsSl ));
    Odrv12 I__4085 (
            .O(N__18125),
            .I(\Lab_UT.sccEmsBitsSl ));
    InMux I__4084 (
            .O(N__18118),
            .I(N__18115));
    LocalMux I__4083 (
            .O(N__18115),
            .I(N__18112));
    Odrv4 I__4082 (
            .O(N__18112),
            .I(\Lab_UT.scctrl.g2 ));
    InMux I__4081 (
            .O(N__18109),
            .I(N__18106));
    LocalMux I__4080 (
            .O(N__18106),
            .I(N__18103));
    Span4Mux_s3_v I__4079 (
            .O(N__18103),
            .I(N__18099));
    InMux I__4078 (
            .O(N__18102),
            .I(N__18096));
    Odrv4 I__4077 (
            .O(N__18099),
            .I(\Lab_UT.scctrl.next_state_rst_3 ));
    LocalMux I__4076 (
            .O(N__18096),
            .I(\Lab_UT.scctrl.next_state_rst_3 ));
    InMux I__4075 (
            .O(N__18091),
            .I(N__18088));
    LocalMux I__4074 (
            .O(N__18088),
            .I(N__18035));
    SRMux I__4073 (
            .O(N__18087),
            .I(N__17932));
    SRMux I__4072 (
            .O(N__18086),
            .I(N__17932));
    SRMux I__4071 (
            .O(N__18085),
            .I(N__17932));
    SRMux I__4070 (
            .O(N__18084),
            .I(N__17932));
    SRMux I__4069 (
            .O(N__18083),
            .I(N__17932));
    SRMux I__4068 (
            .O(N__18082),
            .I(N__17932));
    SRMux I__4067 (
            .O(N__18081),
            .I(N__17932));
    SRMux I__4066 (
            .O(N__18080),
            .I(N__17932));
    SRMux I__4065 (
            .O(N__18079),
            .I(N__17932));
    SRMux I__4064 (
            .O(N__18078),
            .I(N__17932));
    SRMux I__4063 (
            .O(N__18077),
            .I(N__17932));
    SRMux I__4062 (
            .O(N__18076),
            .I(N__17932));
    SRMux I__4061 (
            .O(N__18075),
            .I(N__17932));
    SRMux I__4060 (
            .O(N__18074),
            .I(N__17932));
    SRMux I__4059 (
            .O(N__18073),
            .I(N__17932));
    SRMux I__4058 (
            .O(N__18072),
            .I(N__17932));
    SRMux I__4057 (
            .O(N__18071),
            .I(N__17932));
    SRMux I__4056 (
            .O(N__18070),
            .I(N__17932));
    SRMux I__4055 (
            .O(N__18069),
            .I(N__17932));
    SRMux I__4054 (
            .O(N__18068),
            .I(N__17932));
    SRMux I__4053 (
            .O(N__18067),
            .I(N__17932));
    SRMux I__4052 (
            .O(N__18066),
            .I(N__17932));
    SRMux I__4051 (
            .O(N__18065),
            .I(N__17932));
    SRMux I__4050 (
            .O(N__18064),
            .I(N__17932));
    SRMux I__4049 (
            .O(N__18063),
            .I(N__17932));
    SRMux I__4048 (
            .O(N__18062),
            .I(N__17932));
    SRMux I__4047 (
            .O(N__18061),
            .I(N__17932));
    SRMux I__4046 (
            .O(N__18060),
            .I(N__17932));
    SRMux I__4045 (
            .O(N__18059),
            .I(N__17932));
    SRMux I__4044 (
            .O(N__18058),
            .I(N__17932));
    SRMux I__4043 (
            .O(N__18057),
            .I(N__17932));
    SRMux I__4042 (
            .O(N__18056),
            .I(N__17932));
    SRMux I__4041 (
            .O(N__18055),
            .I(N__17932));
    SRMux I__4040 (
            .O(N__18054),
            .I(N__17932));
    SRMux I__4039 (
            .O(N__18053),
            .I(N__17932));
    SRMux I__4038 (
            .O(N__18052),
            .I(N__17932));
    SRMux I__4037 (
            .O(N__18051),
            .I(N__17932));
    SRMux I__4036 (
            .O(N__18050),
            .I(N__17932));
    SRMux I__4035 (
            .O(N__18049),
            .I(N__17932));
    SRMux I__4034 (
            .O(N__18048),
            .I(N__17932));
    SRMux I__4033 (
            .O(N__18047),
            .I(N__17932));
    SRMux I__4032 (
            .O(N__18046),
            .I(N__17932));
    SRMux I__4031 (
            .O(N__18045),
            .I(N__17932));
    SRMux I__4030 (
            .O(N__18044),
            .I(N__17932));
    SRMux I__4029 (
            .O(N__18043),
            .I(N__17932));
    SRMux I__4028 (
            .O(N__18042),
            .I(N__17932));
    SRMux I__4027 (
            .O(N__18041),
            .I(N__17932));
    SRMux I__4026 (
            .O(N__18040),
            .I(N__17932));
    SRMux I__4025 (
            .O(N__18039),
            .I(N__17932));
    SRMux I__4024 (
            .O(N__18038),
            .I(N__17932));
    Glb2LocalMux I__4023 (
            .O(N__18035),
            .I(N__17932));
    GlobalMux I__4022 (
            .O(N__17932),
            .I(N__17929));
    gio2CtrlBuf I__4021 (
            .O(N__17929),
            .I(resetGen_rst_0_iso_g));
    InMux I__4020 (
            .O(N__17926),
            .I(N__17922));
    InMux I__4019 (
            .O(N__17925),
            .I(N__17919));
    LocalMux I__4018 (
            .O(N__17922),
            .I(N__17916));
    LocalMux I__4017 (
            .O(N__17919),
            .I(N__17913));
    Odrv12 I__4016 (
            .O(N__17916),
            .I(\Lab_UT.scctrl.next_state_rst_2 ));
    Odrv4 I__4015 (
            .O(N__17913),
            .I(\Lab_UT.scctrl.next_state_rst_2 ));
    InMux I__4014 (
            .O(N__17908),
            .I(N__17905));
    LocalMux I__4013 (
            .O(N__17905),
            .I(\Lab_UT.scctrl.N_223_2_reti ));
    InMux I__4012 (
            .O(N__17902),
            .I(N__17899));
    LocalMux I__4011 (
            .O(N__17899),
            .I(N__17894));
    InMux I__4010 (
            .O(N__17898),
            .I(N__17889));
    InMux I__4009 (
            .O(N__17897),
            .I(N__17889));
    Span4Mux_v I__4008 (
            .O(N__17894),
            .I(N__17883));
    LocalMux I__4007 (
            .O(N__17889),
            .I(N__17883));
    InMux I__4006 (
            .O(N__17888),
            .I(N__17879));
    Span4Mux_v I__4005 (
            .O(N__17883),
            .I(N__17876));
    InMux I__4004 (
            .O(N__17882),
            .I(N__17873));
    LocalMux I__4003 (
            .O(N__17879),
            .I(N__17870));
    Odrv4 I__4002 (
            .O(N__17876),
            .I(\Lab_UT.next_state_rst_2_0 ));
    LocalMux I__4001 (
            .O(N__17873),
            .I(\Lab_UT.next_state_rst_2_0 ));
    Odrv4 I__4000 (
            .O(N__17870),
            .I(\Lab_UT.next_state_rst_2_0 ));
    InMux I__3999 (
            .O(N__17863),
            .I(N__17860));
    LocalMux I__3998 (
            .O(N__17860),
            .I(N__17857));
    Span12Mux_s7_v I__3997 (
            .O(N__17857),
            .I(N__17854));
    Odrv12 I__3996 (
            .O(N__17854),
            .I(\Lab_UT.scctrl.g0_i_3 ));
    InMux I__3995 (
            .O(N__17851),
            .I(N__17848));
    LocalMux I__3994 (
            .O(N__17848),
            .I(\Lab_UT.scctrl.N_8 ));
    CascadeMux I__3993 (
            .O(N__17845),
            .I(\Lab_UT.scctrl.g0_i_4_0_cascade_ ));
    InMux I__3992 (
            .O(N__17842),
            .I(N__17833));
    InMux I__3991 (
            .O(N__17841),
            .I(N__17833));
    CascadeMux I__3990 (
            .O(N__17840),
            .I(N__17826));
    InMux I__3989 (
            .O(N__17839),
            .I(N__17821));
    InMux I__3988 (
            .O(N__17838),
            .I(N__17821));
    LocalMux I__3987 (
            .O(N__17833),
            .I(N__17818));
    InMux I__3986 (
            .O(N__17832),
            .I(N__17811));
    InMux I__3985 (
            .O(N__17831),
            .I(N__17811));
    InMux I__3984 (
            .O(N__17830),
            .I(N__17811));
    InMux I__3983 (
            .O(N__17829),
            .I(N__17802));
    InMux I__3982 (
            .O(N__17826),
            .I(N__17802));
    LocalMux I__3981 (
            .O(N__17821),
            .I(N__17799));
    Span4Mux_s3_v I__3980 (
            .O(N__17818),
            .I(N__17794));
    LocalMux I__3979 (
            .O(N__17811),
            .I(N__17794));
    InMux I__3978 (
            .O(N__17810),
            .I(N__17789));
    InMux I__3977 (
            .O(N__17809),
            .I(N__17789));
    IoInMux I__3976 (
            .O(N__17808),
            .I(N__17786));
    IoInMux I__3975 (
            .O(N__17807),
            .I(N__17783));
    LocalMux I__3974 (
            .O(N__17802),
            .I(N__17780));
    Span4Mux_v I__3973 (
            .O(N__17799),
            .I(N__17773));
    Span4Mux_v I__3972 (
            .O(N__17794),
            .I(N__17773));
    LocalMux I__3971 (
            .O(N__17789),
            .I(N__17773));
    LocalMux I__3970 (
            .O(N__17786),
            .I(N__17768));
    LocalMux I__3969 (
            .O(N__17783),
            .I(N__17768));
    Span4Mux_v I__3968 (
            .O(N__17780),
            .I(N__17765));
    Span4Mux_h I__3967 (
            .O(N__17773),
            .I(N__17762));
    Span4Mux_s0_h I__3966 (
            .O(N__17768),
            .I(N__17757));
    Span4Mux_v I__3965 (
            .O(N__17765),
            .I(N__17757));
    Odrv4 I__3964 (
            .O(N__17762),
            .I(led_c_0));
    Odrv4 I__3963 (
            .O(N__17757),
            .I(led_c_0));
    InMux I__3962 (
            .O(N__17752),
            .I(N__17749));
    LocalMux I__3961 (
            .O(N__17749),
            .I(N__17746));
    Odrv4 I__3960 (
            .O(N__17746),
            .I(\Lab_UT.scctrl.N_8_1 ));
    InMux I__3959 (
            .O(N__17743),
            .I(N__17740));
    LocalMux I__3958 (
            .O(N__17740),
            .I(N__17737));
    Odrv4 I__3957 (
            .O(N__17737),
            .I(\Lab_UT.scctrl.N_8_3 ));
    CascadeMux I__3956 (
            .O(N__17734),
            .I(\Lab_UT.scctrl.g0_18_1_cascade_ ));
    InMux I__3955 (
            .O(N__17731),
            .I(N__17727));
    InMux I__3954 (
            .O(N__17730),
            .I(N__17724));
    LocalMux I__3953 (
            .O(N__17727),
            .I(\Lab_UT.scctrl.next_stateZ0Z_2 ));
    LocalMux I__3952 (
            .O(N__17724),
            .I(\Lab_UT.scctrl.next_stateZ0Z_2 ));
    CascadeMux I__3951 (
            .O(N__17719),
            .I(\Lab_UT.scctrl.next_stateZ0Z_2_cascade_ ));
    InMux I__3950 (
            .O(N__17716),
            .I(N__17713));
    LocalMux I__3949 (
            .O(N__17713),
            .I(\Lab_UT.scctrl.N_6_2 ));
    InMux I__3948 (
            .O(N__17710),
            .I(N__17705));
    InMux I__3947 (
            .O(N__17709),
            .I(N__17700));
    InMux I__3946 (
            .O(N__17708),
            .I(N__17700));
    LocalMux I__3945 (
            .O(N__17705),
            .I(\Lab_UT.scctrl.g0_i_3_1 ));
    LocalMux I__3944 (
            .O(N__17700),
            .I(\Lab_UT.scctrl.g0_i_3_1 ));
    CascadeMux I__3943 (
            .O(N__17695),
            .I(N__17692));
    InMux I__3942 (
            .O(N__17692),
            .I(N__17688));
    CascadeMux I__3941 (
            .O(N__17691),
            .I(N__17682));
    LocalMux I__3940 (
            .O(N__17688),
            .I(N__17678));
    InMux I__3939 (
            .O(N__17687),
            .I(N__17675));
    InMux I__3938 (
            .O(N__17686),
            .I(N__17672));
    CascadeMux I__3937 (
            .O(N__17685),
            .I(N__17669));
    InMux I__3936 (
            .O(N__17682),
            .I(N__17666));
    InMux I__3935 (
            .O(N__17681),
            .I(N__17663));
    Span4Mux_s3_v I__3934 (
            .O(N__17678),
            .I(N__17660));
    LocalMux I__3933 (
            .O(N__17675),
            .I(N__17655));
    LocalMux I__3932 (
            .O(N__17672),
            .I(N__17655));
    InMux I__3931 (
            .O(N__17669),
            .I(N__17652));
    LocalMux I__3930 (
            .O(N__17666),
            .I(N__17645));
    LocalMux I__3929 (
            .O(N__17663),
            .I(N__17645));
    Span4Mux_v I__3928 (
            .O(N__17660),
            .I(N__17645));
    Odrv4 I__3927 (
            .O(N__17655),
            .I(next_state_1));
    LocalMux I__3926 (
            .O(N__17652),
            .I(next_state_1));
    Odrv4 I__3925 (
            .O(N__17645),
            .I(next_state_1));
    InMux I__3924 (
            .O(N__17638),
            .I(N__17635));
    LocalMux I__3923 (
            .O(N__17635),
            .I(\Lab_UT.scctrl.g0_i_m4_1_1 ));
    InMux I__3922 (
            .O(N__17632),
            .I(N__17629));
    LocalMux I__3921 (
            .O(N__17629),
            .I(\Lab_UT.scctrl.N_9 ));
    CascadeMux I__3920 (
            .O(N__17626),
            .I(N__17620));
    InMux I__3919 (
            .O(N__17625),
            .I(N__17617));
    CascadeMux I__3918 (
            .O(N__17624),
            .I(N__17612));
    InMux I__3917 (
            .O(N__17623),
            .I(N__17607));
    InMux I__3916 (
            .O(N__17620),
            .I(N__17604));
    LocalMux I__3915 (
            .O(N__17617),
            .I(N__17601));
    InMux I__3914 (
            .O(N__17616),
            .I(N__17598));
    CascadeMux I__3913 (
            .O(N__17615),
            .I(N__17595));
    InMux I__3912 (
            .O(N__17612),
            .I(N__17590));
    InMux I__3911 (
            .O(N__17611),
            .I(N__17590));
    CascadeMux I__3910 (
            .O(N__17610),
            .I(N__17587));
    LocalMux I__3909 (
            .O(N__17607),
            .I(N__17584));
    LocalMux I__3908 (
            .O(N__17604),
            .I(N__17577));
    Span4Mux_h I__3907 (
            .O(N__17601),
            .I(N__17577));
    LocalMux I__3906 (
            .O(N__17598),
            .I(N__17577));
    InMux I__3905 (
            .O(N__17595),
            .I(N__17572));
    LocalMux I__3904 (
            .O(N__17590),
            .I(N__17569));
    InMux I__3903 (
            .O(N__17587),
            .I(N__17566));
    Span4Mux_v I__3902 (
            .O(N__17584),
            .I(N__17561));
    Span4Mux_v I__3901 (
            .O(N__17577),
            .I(N__17561));
    InMux I__3900 (
            .O(N__17576),
            .I(N__17558));
    InMux I__3899 (
            .O(N__17575),
            .I(N__17555));
    LocalMux I__3898 (
            .O(N__17572),
            .I(N__17551));
    Span4Mux_h I__3897 (
            .O(N__17569),
            .I(N__17540));
    LocalMux I__3896 (
            .O(N__17566),
            .I(N__17540));
    Span4Mux_h I__3895 (
            .O(N__17561),
            .I(N__17540));
    LocalMux I__3894 (
            .O(N__17558),
            .I(N__17540));
    LocalMux I__3893 (
            .O(N__17555),
            .I(N__17540));
    InMux I__3892 (
            .O(N__17554),
            .I(N__17537));
    Span4Mux_h I__3891 (
            .O(N__17551),
            .I(N__17534));
    Span4Mux_v I__3890 (
            .O(N__17540),
            .I(N__17531));
    LocalMux I__3889 (
            .O(N__17537),
            .I(rst_i_3_rep2));
    Odrv4 I__3888 (
            .O(N__17534),
            .I(rst_i_3_rep2));
    Odrv4 I__3887 (
            .O(N__17531),
            .I(rst_i_3_rep2));
    InMux I__3886 (
            .O(N__17524),
            .I(N__17521));
    LocalMux I__3885 (
            .O(N__17521),
            .I(N__17517));
    InMux I__3884 (
            .O(N__17520),
            .I(N__17514));
    Odrv4 I__3883 (
            .O(N__17517),
            .I(\Lab_UT.state_ret_8_rep1_RNIJDTUE_1 ));
    LocalMux I__3882 (
            .O(N__17514),
            .I(\Lab_UT.state_ret_8_rep1_RNIJDTUE_1 ));
    CascadeMux I__3881 (
            .O(N__17509),
            .I(\Lab_UT.scctrl.next_state_rst_0_5_0_cascade_ ));
    CascadeMux I__3880 (
            .O(N__17506),
            .I(N__17503));
    InMux I__3879 (
            .O(N__17503),
            .I(N__17491));
    InMux I__3878 (
            .O(N__17502),
            .I(N__17486));
    InMux I__3877 (
            .O(N__17501),
            .I(N__17483));
    InMux I__3876 (
            .O(N__17500),
            .I(N__17477));
    InMux I__3875 (
            .O(N__17499),
            .I(N__17477));
    InMux I__3874 (
            .O(N__17498),
            .I(N__17472));
    InMux I__3873 (
            .O(N__17497),
            .I(N__17469));
    InMux I__3872 (
            .O(N__17496),
            .I(N__17464));
    InMux I__3871 (
            .O(N__17495),
            .I(N__17464));
    InMux I__3870 (
            .O(N__17494),
            .I(N__17461));
    LocalMux I__3869 (
            .O(N__17491),
            .I(N__17458));
    InMux I__3868 (
            .O(N__17490),
            .I(N__17453));
    InMux I__3867 (
            .O(N__17489),
            .I(N__17453));
    LocalMux I__3866 (
            .O(N__17486),
            .I(N__17450));
    LocalMux I__3865 (
            .O(N__17483),
            .I(N__17447));
    InMux I__3864 (
            .O(N__17482),
            .I(N__17443));
    LocalMux I__3863 (
            .O(N__17477),
            .I(N__17437));
    InMux I__3862 (
            .O(N__17476),
            .I(N__17432));
    InMux I__3861 (
            .O(N__17475),
            .I(N__17432));
    LocalMux I__3860 (
            .O(N__17472),
            .I(N__17429));
    LocalMux I__3859 (
            .O(N__17469),
            .I(N__17426));
    LocalMux I__3858 (
            .O(N__17464),
            .I(N__17417));
    LocalMux I__3857 (
            .O(N__17461),
            .I(N__17417));
    Span4Mux_s3_h I__3856 (
            .O(N__17458),
            .I(N__17417));
    LocalMux I__3855 (
            .O(N__17453),
            .I(N__17417));
    Span4Mux_h I__3854 (
            .O(N__17450),
            .I(N__17412));
    Span4Mux_v I__3853 (
            .O(N__17447),
            .I(N__17412));
    InMux I__3852 (
            .O(N__17446),
            .I(N__17409));
    LocalMux I__3851 (
            .O(N__17443),
            .I(N__17406));
    InMux I__3850 (
            .O(N__17442),
            .I(N__17401));
    InMux I__3849 (
            .O(N__17441),
            .I(N__17401));
    InMux I__3848 (
            .O(N__17440),
            .I(N__17398));
    Span4Mux_h I__3847 (
            .O(N__17437),
            .I(N__17393));
    LocalMux I__3846 (
            .O(N__17432),
            .I(N__17393));
    Span12Mux_s4_v I__3845 (
            .O(N__17429),
            .I(N__17388));
    Span12Mux_s11_v I__3844 (
            .O(N__17426),
            .I(N__17388));
    Span4Mux_v I__3843 (
            .O(N__17417),
            .I(N__17383));
    Span4Mux_v I__3842 (
            .O(N__17412),
            .I(N__17383));
    LocalMux I__3841 (
            .O(N__17409),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    Odrv12 I__3840 (
            .O(N__17406),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    LocalMux I__3839 (
            .O(N__17401),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    LocalMux I__3838 (
            .O(N__17398),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    Odrv4 I__3837 (
            .O(N__17393),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    Odrv12 I__3836 (
            .O(N__17388),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    Odrv4 I__3835 (
            .O(N__17383),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    CascadeMux I__3834 (
            .O(N__17368),
            .I(N__17364));
    InMux I__3833 (
            .O(N__17367),
            .I(N__17360));
    InMux I__3832 (
            .O(N__17364),
            .I(N__17356));
    InMux I__3831 (
            .O(N__17363),
            .I(N__17353));
    LocalMux I__3830 (
            .O(N__17360),
            .I(N__17350));
    InMux I__3829 (
            .O(N__17359),
            .I(N__17347));
    LocalMux I__3828 (
            .O(N__17356),
            .I(N__17344));
    LocalMux I__3827 (
            .O(N__17353),
            .I(N__17340));
    Span4Mux_v I__3826 (
            .O(N__17350),
            .I(N__17337));
    LocalMux I__3825 (
            .O(N__17347),
            .I(N__17333));
    Span4Mux_h I__3824 (
            .O(N__17344),
            .I(N__17330));
    InMux I__3823 (
            .O(N__17343),
            .I(N__17327));
    Span4Mux_h I__3822 (
            .O(N__17340),
            .I(N__17324));
    Span4Mux_v I__3821 (
            .O(N__17337),
            .I(N__17321));
    InMux I__3820 (
            .O(N__17336),
            .I(N__17318));
    Span4Mux_h I__3819 (
            .O(N__17333),
            .I(N__17315));
    Sp12to4 I__3818 (
            .O(N__17330),
            .I(N__17310));
    LocalMux I__3817 (
            .O(N__17327),
            .I(N__17310));
    Odrv4 I__3816 (
            .O(N__17324),
            .I(rst_i_3_rep1));
    Odrv4 I__3815 (
            .O(N__17321),
            .I(rst_i_3_rep1));
    LocalMux I__3814 (
            .O(N__17318),
            .I(rst_i_3_rep1));
    Odrv4 I__3813 (
            .O(N__17315),
            .I(rst_i_3_rep1));
    Odrv12 I__3812 (
            .O(N__17310),
            .I(rst_i_3_rep1));
    InMux I__3811 (
            .O(N__17299),
            .I(N__17296));
    LocalMux I__3810 (
            .O(N__17296),
            .I(\Lab_UT.scctrl.g0_i_a8_1 ));
    CascadeMux I__3809 (
            .O(N__17293),
            .I(N__17290));
    InMux I__3808 (
            .O(N__17290),
            .I(N__17287));
    LocalMux I__3807 (
            .O(N__17287),
            .I(\Lab_UT.scctrl.g0_i_0_0 ));
    InMux I__3806 (
            .O(N__17284),
            .I(N__17281));
    LocalMux I__3805 (
            .O(N__17281),
            .I(N__17278));
    Odrv4 I__3804 (
            .O(N__17278),
            .I(\Lab_UT.scctrl.g0_7_3 ));
    CascadeMux I__3803 (
            .O(N__17275),
            .I(N__17272));
    InMux I__3802 (
            .O(N__17272),
            .I(N__17269));
    LocalMux I__3801 (
            .O(N__17269),
            .I(\Lab_UT.scctrl.g0_7_2 ));
    CascadeMux I__3800 (
            .O(N__17266),
            .I(\Lab_UT.scctrl.g2_cascade_ ));
    InMux I__3799 (
            .O(N__17263),
            .I(N__17260));
    LocalMux I__3798 (
            .O(N__17260),
            .I(\Lab_UT.scctrl.g1_1 ));
    InMux I__3797 (
            .O(N__17257),
            .I(N__17254));
    LocalMux I__3796 (
            .O(N__17254),
            .I(N__17251));
    Odrv4 I__3795 (
            .O(N__17251),
            .I(\Lab_UT.scctrl.g0_1_0 ));
    CascadeMux I__3794 (
            .O(N__17248),
            .I(\Lab_UT.scctrl.N_222i_cascade_ ));
    InMux I__3793 (
            .O(N__17245),
            .I(N__17242));
    LocalMux I__3792 (
            .O(N__17242),
            .I(\Lab_UT.scctrl.N_223_1_reti ));
    InMux I__3791 (
            .O(N__17239),
            .I(N__17236));
    LocalMux I__3790 (
            .O(N__17236),
            .I(N__17233));
    Span4Mux_h I__3789 (
            .O(N__17233),
            .I(N__17230));
    Odrv4 I__3788 (
            .O(N__17230),
            .I(shifter_0_fast_RNI639J4_2));
    CascadeMux I__3787 (
            .O(N__17227),
            .I(\Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433_cascade_ ));
    InMux I__3786 (
            .O(N__17224),
            .I(N__17221));
    LocalMux I__3785 (
            .O(N__17221),
            .I(\Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0 ));
    InMux I__3784 (
            .O(N__17218),
            .I(N__17212));
    InMux I__3783 (
            .O(N__17217),
            .I(N__17205));
    InMux I__3782 (
            .O(N__17216),
            .I(N__17205));
    InMux I__3781 (
            .O(N__17215),
            .I(N__17205));
    LocalMux I__3780 (
            .O(N__17212),
            .I(N__17202));
    LocalMux I__3779 (
            .O(N__17205),
            .I(N__17199));
    Span4Mux_v I__3778 (
            .O(N__17202),
            .I(N__17195));
    Span4Mux_h I__3777 (
            .O(N__17199),
            .I(N__17192));
    InMux I__3776 (
            .O(N__17198),
            .I(N__17189));
    Odrv4 I__3775 (
            .O(N__17195),
            .I(\Lab_UT.de_bigD ));
    Odrv4 I__3774 (
            .O(N__17192),
            .I(\Lab_UT.de_bigD ));
    LocalMux I__3773 (
            .O(N__17189),
            .I(\Lab_UT.de_bigD ));
    InMux I__3772 (
            .O(N__17182),
            .I(N__17179));
    LocalMux I__3771 (
            .O(N__17179),
            .I(N__17175));
    CascadeMux I__3770 (
            .O(N__17178),
            .I(N__17171));
    Span4Mux_v I__3769 (
            .O(N__17175),
            .I(N__17167));
    InMux I__3768 (
            .O(N__17174),
            .I(N__17160));
    InMux I__3767 (
            .O(N__17171),
            .I(N__17160));
    InMux I__3766 (
            .O(N__17170),
            .I(N__17160));
    Odrv4 I__3765 (
            .O(N__17167),
            .I(\Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433 ));
    LocalMux I__3764 (
            .O(N__17160),
            .I(\Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433 ));
    CascadeMux I__3763 (
            .O(N__17155),
            .I(N__17151));
    InMux I__3762 (
            .O(N__17154),
            .I(N__17145));
    InMux I__3761 (
            .O(N__17151),
            .I(N__17136));
    InMux I__3760 (
            .O(N__17150),
            .I(N__17136));
    InMux I__3759 (
            .O(N__17149),
            .I(N__17136));
    InMux I__3758 (
            .O(N__17148),
            .I(N__17136));
    LocalMux I__3757 (
            .O(N__17145),
            .I(N__17132));
    LocalMux I__3756 (
            .O(N__17136),
            .I(N__17129));
    InMux I__3755 (
            .O(N__17135),
            .I(N__17126));
    Odrv4 I__3754 (
            .O(N__17132),
            .I(\Lab_UT.de_bigL ));
    Odrv12 I__3753 (
            .O(N__17129),
            .I(\Lab_UT.de_bigL ));
    LocalMux I__3752 (
            .O(N__17126),
            .I(\Lab_UT.de_bigL ));
    CascadeMux I__3751 (
            .O(N__17119),
            .I(N__17116));
    InMux I__3750 (
            .O(N__17116),
            .I(N__17113));
    LocalMux I__3749 (
            .O(N__17113),
            .I(N__17107));
    InMux I__3748 (
            .O(N__17112),
            .I(N__17100));
    InMux I__3747 (
            .O(N__17111),
            .I(N__17100));
    InMux I__3746 (
            .O(N__17110),
            .I(N__17100));
    Odrv4 I__3745 (
            .O(N__17107),
            .I(\Lab_UT.scctrl.next_state_1_i_o2_0_d_1 ));
    LocalMux I__3744 (
            .O(N__17100),
            .I(\Lab_UT.scctrl.next_state_1_i_o2_0_d_1 ));
    CascadeMux I__3743 (
            .O(N__17095),
            .I(N__17092));
    InMux I__3742 (
            .O(N__17092),
            .I(N__17086));
    InMux I__3741 (
            .O(N__17091),
            .I(N__17086));
    LocalMux I__3740 (
            .O(N__17086),
            .I(N__17083));
    Span4Mux_v I__3739 (
            .O(N__17083),
            .I(N__17080));
    Odrv4 I__3738 (
            .O(N__17080),
            .I(\Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0Z_2 ));
    InMux I__3737 (
            .O(N__17077),
            .I(N__17067));
    InMux I__3736 (
            .O(N__17076),
            .I(N__17067));
    InMux I__3735 (
            .O(N__17075),
            .I(N__17063));
    InMux I__3734 (
            .O(N__17074),
            .I(N__17060));
    InMux I__3733 (
            .O(N__17073),
            .I(N__17056));
    InMux I__3732 (
            .O(N__17072),
            .I(N__17053));
    LocalMux I__3731 (
            .O(N__17067),
            .I(N__17050));
    InMux I__3730 (
            .O(N__17066),
            .I(N__17045));
    LocalMux I__3729 (
            .O(N__17063),
            .I(N__17042));
    LocalMux I__3728 (
            .O(N__17060),
            .I(N__17039));
    InMux I__3727 (
            .O(N__17059),
            .I(N__17036));
    LocalMux I__3726 (
            .O(N__17056),
            .I(N__17031));
    LocalMux I__3725 (
            .O(N__17053),
            .I(N__17031));
    Span4Mux_v I__3724 (
            .O(N__17050),
            .I(N__17028));
    InMux I__3723 (
            .O(N__17049),
            .I(N__17023));
    InMux I__3722 (
            .O(N__17048),
            .I(N__17023));
    LocalMux I__3721 (
            .O(N__17045),
            .I(N__17016));
    Span4Mux_h I__3720 (
            .O(N__17042),
            .I(N__17011));
    Span4Mux_h I__3719 (
            .O(N__17039),
            .I(N__17011));
    LocalMux I__3718 (
            .O(N__17036),
            .I(N__17008));
    Span4Mux_h I__3717 (
            .O(N__17031),
            .I(N__17005));
    Span4Mux_s3_h I__3716 (
            .O(N__17028),
            .I(N__17002));
    LocalMux I__3715 (
            .O(N__17023),
            .I(N__16999));
    InMux I__3714 (
            .O(N__17022),
            .I(N__16994));
    InMux I__3713 (
            .O(N__17021),
            .I(N__16994));
    InMux I__3712 (
            .O(N__17020),
            .I(N__16989));
    InMux I__3711 (
            .O(N__17019),
            .I(N__16989));
    Odrv4 I__3710 (
            .O(N__17016),
            .I(bu_rx_data_6));
    Odrv4 I__3709 (
            .O(N__17011),
            .I(bu_rx_data_6));
    Odrv4 I__3708 (
            .O(N__17008),
            .I(bu_rx_data_6));
    Odrv4 I__3707 (
            .O(N__17005),
            .I(bu_rx_data_6));
    Odrv4 I__3706 (
            .O(N__17002),
            .I(bu_rx_data_6));
    Odrv4 I__3705 (
            .O(N__16999),
            .I(bu_rx_data_6));
    LocalMux I__3704 (
            .O(N__16994),
            .I(bu_rx_data_6));
    LocalMux I__3703 (
            .O(N__16989),
            .I(bu_rx_data_6));
    CascadeMux I__3702 (
            .O(N__16972),
            .I(N__16967));
    CascadeMux I__3701 (
            .O(N__16971),
            .I(N__16961));
    InMux I__3700 (
            .O(N__16970),
            .I(N__16951));
    InMux I__3699 (
            .O(N__16967),
            .I(N__16946));
    InMux I__3698 (
            .O(N__16966),
            .I(N__16946));
    InMux I__3697 (
            .O(N__16965),
            .I(N__16937));
    InMux I__3696 (
            .O(N__16964),
            .I(N__16934));
    InMux I__3695 (
            .O(N__16961),
            .I(N__16931));
    InMux I__3694 (
            .O(N__16960),
            .I(N__16928));
    InMux I__3693 (
            .O(N__16959),
            .I(N__16921));
    InMux I__3692 (
            .O(N__16958),
            .I(N__16921));
    InMux I__3691 (
            .O(N__16957),
            .I(N__16921));
    InMux I__3690 (
            .O(N__16956),
            .I(N__16918));
    InMux I__3689 (
            .O(N__16955),
            .I(N__16915));
    InMux I__3688 (
            .O(N__16954),
            .I(N__16912));
    LocalMux I__3687 (
            .O(N__16951),
            .I(N__16909));
    LocalMux I__3686 (
            .O(N__16946),
            .I(N__16906));
    InMux I__3685 (
            .O(N__16945),
            .I(N__16901));
    InMux I__3684 (
            .O(N__16944),
            .I(N__16901));
    InMux I__3683 (
            .O(N__16943),
            .I(N__16896));
    InMux I__3682 (
            .O(N__16942),
            .I(N__16891));
    InMux I__3681 (
            .O(N__16941),
            .I(N__16891));
    CascadeMux I__3680 (
            .O(N__16940),
            .I(N__16887));
    LocalMux I__3679 (
            .O(N__16937),
            .I(N__16883));
    LocalMux I__3678 (
            .O(N__16934),
            .I(N__16880));
    LocalMux I__3677 (
            .O(N__16931),
            .I(N__16874));
    LocalMux I__3676 (
            .O(N__16928),
            .I(N__16867));
    LocalMux I__3675 (
            .O(N__16921),
            .I(N__16867));
    LocalMux I__3674 (
            .O(N__16918),
            .I(N__16867));
    LocalMux I__3673 (
            .O(N__16915),
            .I(N__16864));
    LocalMux I__3672 (
            .O(N__16912),
            .I(N__16855));
    Span4Mux_v I__3671 (
            .O(N__16909),
            .I(N__16855));
    Span4Mux_v I__3670 (
            .O(N__16906),
            .I(N__16855));
    LocalMux I__3669 (
            .O(N__16901),
            .I(N__16855));
    CascadeMux I__3668 (
            .O(N__16900),
            .I(N__16850));
    CascadeMux I__3667 (
            .O(N__16899),
            .I(N__16847));
    LocalMux I__3666 (
            .O(N__16896),
            .I(N__16843));
    LocalMux I__3665 (
            .O(N__16891),
            .I(N__16840));
    InMux I__3664 (
            .O(N__16890),
            .I(N__16833));
    InMux I__3663 (
            .O(N__16887),
            .I(N__16833));
    InMux I__3662 (
            .O(N__16886),
            .I(N__16833));
    Span4Mux_h I__3661 (
            .O(N__16883),
            .I(N__16828));
    Span4Mux_h I__3660 (
            .O(N__16880),
            .I(N__16828));
    InMux I__3659 (
            .O(N__16879),
            .I(N__16825));
    InMux I__3658 (
            .O(N__16878),
            .I(N__16820));
    InMux I__3657 (
            .O(N__16877),
            .I(N__16820));
    Span4Mux_v I__3656 (
            .O(N__16874),
            .I(N__16815));
    Span4Mux_v I__3655 (
            .O(N__16867),
            .I(N__16815));
    Span4Mux_h I__3654 (
            .O(N__16864),
            .I(N__16810));
    Span4Mux_h I__3653 (
            .O(N__16855),
            .I(N__16810));
    InMux I__3652 (
            .O(N__16854),
            .I(N__16801));
    InMux I__3651 (
            .O(N__16853),
            .I(N__16801));
    InMux I__3650 (
            .O(N__16850),
            .I(N__16801));
    InMux I__3649 (
            .O(N__16847),
            .I(N__16801));
    InMux I__3648 (
            .O(N__16846),
            .I(N__16798));
    Span4Mux_v I__3647 (
            .O(N__16843),
            .I(N__16791));
    Span4Mux_v I__3646 (
            .O(N__16840),
            .I(N__16791));
    LocalMux I__3645 (
            .O(N__16833),
            .I(N__16791));
    Odrv4 I__3644 (
            .O(N__16828),
            .I(bu_rx_data_7));
    LocalMux I__3643 (
            .O(N__16825),
            .I(bu_rx_data_7));
    LocalMux I__3642 (
            .O(N__16820),
            .I(bu_rx_data_7));
    Odrv4 I__3641 (
            .O(N__16815),
            .I(bu_rx_data_7));
    Odrv4 I__3640 (
            .O(N__16810),
            .I(bu_rx_data_7));
    LocalMux I__3639 (
            .O(N__16801),
            .I(bu_rx_data_7));
    LocalMux I__3638 (
            .O(N__16798),
            .I(bu_rx_data_7));
    Odrv4 I__3637 (
            .O(N__16791),
            .I(bu_rx_data_7));
    InMux I__3636 (
            .O(N__16774),
            .I(N__16771));
    LocalMux I__3635 (
            .O(N__16771),
            .I(N__16768));
    Span4Mux_v I__3634 (
            .O(N__16768),
            .I(N__16765));
    Sp12to4 I__3633 (
            .O(N__16765),
            .I(N__16762));
    Odrv12 I__3632 (
            .O(N__16762),
            .I(resetGen_escKey_4));
    CEMux I__3631 (
            .O(N__16759),
            .I(N__16735));
    CEMux I__3630 (
            .O(N__16758),
            .I(N__16735));
    CEMux I__3629 (
            .O(N__16757),
            .I(N__16735));
    CEMux I__3628 (
            .O(N__16756),
            .I(N__16735));
    CEMux I__3627 (
            .O(N__16755),
            .I(N__16735));
    CEMux I__3626 (
            .O(N__16754),
            .I(N__16735));
    CEMux I__3625 (
            .O(N__16753),
            .I(N__16735));
    CEMux I__3624 (
            .O(N__16752),
            .I(N__16735));
    GlobalMux I__3623 (
            .O(N__16735),
            .I(N__16732));
    gio2CtrlBuf I__3622 (
            .O(N__16732),
            .I(N_41_i_g));
    InMux I__3621 (
            .O(N__16729),
            .I(N__16726));
    LocalMux I__3620 (
            .O(N__16726),
            .I(N__16723));
    Span4Mux_v I__3619 (
            .O(N__16723),
            .I(N__16720));
    Span4Mux_s2_h I__3618 (
            .O(N__16720),
            .I(N__16717));
    Span4Mux_h I__3617 (
            .O(N__16717),
            .I(N__16714));
    Odrv4 I__3616 (
            .O(N__16714),
            .I(\Lab_UT.scctrl.g0_2_1 ));
    InMux I__3615 (
            .O(N__16711),
            .I(N__16708));
    LocalMux I__3614 (
            .O(N__16708),
            .I(\Lab_UT.scctrl.next_state_rst_0_3_N_6_0 ));
    CascadeMux I__3613 (
            .O(N__16705),
            .I(\Lab_UT.scctrl.g1_0_0_cascade_ ));
    InMux I__3612 (
            .O(N__16702),
            .I(N__16699));
    LocalMux I__3611 (
            .O(N__16699),
            .I(N__16696));
    Odrv12 I__3610 (
            .O(N__16696),
            .I(\Lab_UT.scctrl.g0_1_3 ));
    InMux I__3609 (
            .O(N__16693),
            .I(N__16690));
    LocalMux I__3608 (
            .O(N__16690),
            .I(N__16687));
    Odrv4 I__3607 (
            .O(N__16687),
            .I(\Lab_UT.scctrl.g0_1_0_0 ));
    CascadeMux I__3606 (
            .O(N__16684),
            .I(\Lab_UT.scctrl.N_127_i_i_o6_0_1_cascade_ ));
    InMux I__3605 (
            .O(N__16681),
            .I(N__16678));
    LocalMux I__3604 (
            .O(N__16678),
            .I(\Lab_UT.scctrl.N_127_i_i_a6_1 ));
    InMux I__3603 (
            .O(N__16675),
            .I(N__16672));
    LocalMux I__3602 (
            .O(N__16672),
            .I(\Lab_UT.scctrl.N_190_0_0 ));
    InMux I__3601 (
            .O(N__16669),
            .I(N__16664));
    InMux I__3600 (
            .O(N__16668),
            .I(N__16659));
    InMux I__3599 (
            .O(N__16667),
            .I(N__16659));
    LocalMux I__3598 (
            .O(N__16664),
            .I(N__16656));
    LocalMux I__3597 (
            .O(N__16659),
            .I(N__16653));
    Span4Mux_h I__3596 (
            .O(N__16656),
            .I(N__16650));
    Span4Mux_s3_h I__3595 (
            .O(N__16653),
            .I(N__16647));
    Odrv4 I__3594 (
            .O(N__16650),
            .I(\Lab_UT.next_state_rst_0_5 ));
    Odrv4 I__3593 (
            .O(N__16647),
            .I(\Lab_UT.next_state_rst_0_5 ));
    InMux I__3592 (
            .O(N__16642),
            .I(N__16639));
    LocalMux I__3591 (
            .O(N__16639),
            .I(\Lab_UT.scdp.a2b.N_6_4 ));
    CascadeMux I__3590 (
            .O(N__16636),
            .I(N__16633));
    InMux I__3589 (
            .O(N__16633),
            .I(N__16630));
    LocalMux I__3588 (
            .O(N__16630),
            .I(N__16627));
    Odrv4 I__3587 (
            .O(N__16627),
            .I(\Lab_UT.state_ret_8_rep1_RNIHA8U3 ));
    InMux I__3586 (
            .O(N__16624),
            .I(N__16618));
    InMux I__3585 (
            .O(N__16623),
            .I(N__16618));
    LocalMux I__3584 (
            .O(N__16618),
            .I(\Lab_UT.N_182 ));
    InMux I__3583 (
            .O(N__16615),
            .I(N__16612));
    LocalMux I__3582 (
            .O(N__16612),
            .I(\Lab_UT.scdp.a2b.g0_iZ0Z_9 ));
    InMux I__3581 (
            .O(N__16609),
            .I(N__16606));
    LocalMux I__3580 (
            .O(N__16606),
            .I(N__16600));
    InMux I__3579 (
            .O(N__16605),
            .I(N__16593));
    InMux I__3578 (
            .O(N__16604),
            .I(N__16593));
    InMux I__3577 (
            .O(N__16603),
            .I(N__16593));
    Odrv4 I__3576 (
            .O(N__16600),
            .I(\Lab_UT.state_2_RNI3PVB9_2 ));
    LocalMux I__3575 (
            .O(N__16593),
            .I(\Lab_UT.state_2_RNI3PVB9_2 ));
    InMux I__3574 (
            .O(N__16588),
            .I(N__16585));
    LocalMux I__3573 (
            .O(N__16585),
            .I(\Lab_UT.scctrl.N_182_0 ));
    CascadeMux I__3572 (
            .O(N__16582),
            .I(N__16578));
    InMux I__3571 (
            .O(N__16581),
            .I(N__16575));
    InMux I__3570 (
            .O(N__16578),
            .I(N__16572));
    LocalMux I__3569 (
            .O(N__16575),
            .I(N__16569));
    LocalMux I__3568 (
            .O(N__16572),
            .I(N__16566));
    Odrv12 I__3567 (
            .O(N__16569),
            .I(\Lab_UT.scctrl.N_166_0_1 ));
    Odrv4 I__3566 (
            .O(N__16566),
            .I(\Lab_UT.scctrl.N_166_0_1 ));
    InMux I__3565 (
            .O(N__16561),
            .I(N__16557));
    InMux I__3564 (
            .O(N__16560),
            .I(N__16554));
    LocalMux I__3563 (
            .O(N__16557),
            .I(N__16551));
    LocalMux I__3562 (
            .O(N__16554),
            .I(N__16541));
    Span4Mux_v I__3561 (
            .O(N__16551),
            .I(N__16541));
    InMux I__3560 (
            .O(N__16550),
            .I(N__16538));
    InMux I__3559 (
            .O(N__16549),
            .I(N__16535));
    InMux I__3558 (
            .O(N__16548),
            .I(N__16532));
    InMux I__3557 (
            .O(N__16547),
            .I(N__16527));
    InMux I__3556 (
            .O(N__16546),
            .I(N__16527));
    Span4Mux_h I__3555 (
            .O(N__16541),
            .I(N__16520));
    LocalMux I__3554 (
            .O(N__16538),
            .I(N__16520));
    LocalMux I__3553 (
            .O(N__16535),
            .I(N__16520));
    LocalMux I__3552 (
            .O(N__16532),
            .I(bu_rx_data_0_rep1));
    LocalMux I__3551 (
            .O(N__16527),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__3550 (
            .O(N__16520),
            .I(bu_rx_data_0_rep1));
    CascadeMux I__3549 (
            .O(N__16513),
            .I(\Lab_UT.scctrl.next_state_1_i_o2_0_d_1_cascade_ ));
    InMux I__3548 (
            .O(N__16510),
            .I(N__16506));
    InMux I__3547 (
            .O(N__16509),
            .I(N__16501));
    LocalMux I__3546 (
            .O(N__16506),
            .I(N__16497));
    CascadeMux I__3545 (
            .O(N__16505),
            .I(N__16494));
    CascadeMux I__3544 (
            .O(N__16504),
            .I(N__16491));
    LocalMux I__3543 (
            .O(N__16501),
            .I(N__16486));
    InMux I__3542 (
            .O(N__16500),
            .I(N__16483));
    Span4Mux_h I__3541 (
            .O(N__16497),
            .I(N__16480));
    InMux I__3540 (
            .O(N__16494),
            .I(N__16477));
    InMux I__3539 (
            .O(N__16491),
            .I(N__16474));
    InMux I__3538 (
            .O(N__16490),
            .I(N__16471));
    InMux I__3537 (
            .O(N__16489),
            .I(N__16468));
    Span4Mux_h I__3536 (
            .O(N__16486),
            .I(N__16463));
    LocalMux I__3535 (
            .O(N__16483),
            .I(N__16463));
    Odrv4 I__3534 (
            .O(N__16480),
            .I(buart__rx_shifter_0_fast_2));
    LocalMux I__3533 (
            .O(N__16477),
            .I(buart__rx_shifter_0_fast_2));
    LocalMux I__3532 (
            .O(N__16474),
            .I(buart__rx_shifter_0_fast_2));
    LocalMux I__3531 (
            .O(N__16471),
            .I(buart__rx_shifter_0_fast_2));
    LocalMux I__3530 (
            .O(N__16468),
            .I(buart__rx_shifter_0_fast_2));
    Odrv4 I__3529 (
            .O(N__16463),
            .I(buart__rx_shifter_0_fast_2));
    CascadeMux I__3528 (
            .O(N__16450),
            .I(\Lab_UT.scctrl.next_state_rst_0_3_N_5L8Z0Z_1_cascade_ ));
    InMux I__3527 (
            .O(N__16447),
            .I(N__16443));
    InMux I__3526 (
            .O(N__16446),
            .I(N__16440));
    LocalMux I__3525 (
            .O(N__16443),
            .I(N__16437));
    LocalMux I__3524 (
            .O(N__16440),
            .I(N__16434));
    Span4Mux_v I__3523 (
            .O(N__16437),
            .I(N__16427));
    Span4Mux_h I__3522 (
            .O(N__16434),
            .I(N__16427));
    InMux I__3521 (
            .O(N__16433),
            .I(N__16422));
    InMux I__3520 (
            .O(N__16432),
            .I(N__16422));
    Odrv4 I__3519 (
            .O(N__16427),
            .I(Lab_UT_dk_de_bigD_6));
    LocalMux I__3518 (
            .O(N__16422),
            .I(Lab_UT_dk_de_bigD_6));
    CascadeMux I__3517 (
            .O(N__16417),
            .I(N__16414));
    InMux I__3516 (
            .O(N__16414),
            .I(N__16411));
    LocalMux I__3515 (
            .O(N__16411),
            .I(\Lab_UT.scctrl.g0_0_i_1_1 ));
    CascadeMux I__3514 (
            .O(N__16408),
            .I(N__16405));
    InMux I__3513 (
            .O(N__16405),
            .I(N__16402));
    LocalMux I__3512 (
            .O(N__16402),
            .I(N__16399));
    Span4Mux_h I__3511 (
            .O(N__16399),
            .I(N__16396));
    Odrv4 I__3510 (
            .O(N__16396),
            .I(\Lab_UT.scctrl.N_14 ));
    InMux I__3509 (
            .O(N__16393),
            .I(N__16390));
    LocalMux I__3508 (
            .O(N__16390),
            .I(\Lab_UT.scdp.a2b.g0_iZ0Z_4 ));
    InMux I__3507 (
            .O(N__16387),
            .I(N__16384));
    LocalMux I__3506 (
            .O(N__16384),
            .I(\Lab_UT.N_5 ));
    CascadeMux I__3505 (
            .O(N__16381),
            .I(\Lab_UT.scdp.a2b.g0_iZ0Z_8_cascade_ ));
    InMux I__3504 (
            .O(N__16378),
            .I(N__16375));
    LocalMux I__3503 (
            .O(N__16375),
            .I(\Lab_UT.scdp.a2b.g0_3_a3_6 ));
    CascadeMux I__3502 (
            .O(N__16372),
            .I(N__16368));
    InMux I__3501 (
            .O(N__16371),
            .I(N__16364));
    InMux I__3500 (
            .O(N__16368),
            .I(N__16359));
    InMux I__3499 (
            .O(N__16367),
            .I(N__16359));
    LocalMux I__3498 (
            .O(N__16364),
            .I(N__16355));
    LocalMux I__3497 (
            .O(N__16359),
            .I(N__16349));
    InMux I__3496 (
            .O(N__16358),
            .I(N__16346));
    Span4Mux_v I__3495 (
            .O(N__16355),
            .I(N__16343));
    InMux I__3494 (
            .O(N__16354),
            .I(N__16338));
    InMux I__3493 (
            .O(N__16353),
            .I(N__16333));
    InMux I__3492 (
            .O(N__16352),
            .I(N__16333));
    Span4Mux_v I__3491 (
            .O(N__16349),
            .I(N__16330));
    LocalMux I__3490 (
            .O(N__16346),
            .I(N__16327));
    Span4Mux_s2_h I__3489 (
            .O(N__16343),
            .I(N__16324));
    InMux I__3488 (
            .O(N__16342),
            .I(N__16319));
    InMux I__3487 (
            .O(N__16341),
            .I(N__16319));
    LocalMux I__3486 (
            .O(N__16338),
            .I(\Lab_UT.de_cr_2 ));
    LocalMux I__3485 (
            .O(N__16333),
            .I(\Lab_UT.de_cr_2 ));
    Odrv4 I__3484 (
            .O(N__16330),
            .I(\Lab_UT.de_cr_2 ));
    Odrv4 I__3483 (
            .O(N__16327),
            .I(\Lab_UT.de_cr_2 ));
    Odrv4 I__3482 (
            .O(N__16324),
            .I(\Lab_UT.de_cr_2 ));
    LocalMux I__3481 (
            .O(N__16319),
            .I(\Lab_UT.de_cr_2 ));
    InMux I__3480 (
            .O(N__16306),
            .I(N__16301));
    InMux I__3479 (
            .O(N__16305),
            .I(N__16298));
    CascadeMux I__3478 (
            .O(N__16304),
            .I(N__16294));
    LocalMux I__3477 (
            .O(N__16301),
            .I(N__16286));
    LocalMux I__3476 (
            .O(N__16298),
            .I(N__16286));
    InMux I__3475 (
            .O(N__16297),
            .I(N__16283));
    InMux I__3474 (
            .O(N__16294),
            .I(N__16280));
    CascadeMux I__3473 (
            .O(N__16293),
            .I(N__16277));
    CascadeMux I__3472 (
            .O(N__16292),
            .I(N__16274));
    CascadeMux I__3471 (
            .O(N__16291),
            .I(N__16271));
    Span4Mux_v I__3470 (
            .O(N__16286),
            .I(N__16267));
    LocalMux I__3469 (
            .O(N__16283),
            .I(N__16264));
    LocalMux I__3468 (
            .O(N__16280),
            .I(N__16261));
    InMux I__3467 (
            .O(N__16277),
            .I(N__16256));
    InMux I__3466 (
            .O(N__16274),
            .I(N__16256));
    InMux I__3465 (
            .O(N__16271),
            .I(N__16251));
    InMux I__3464 (
            .O(N__16270),
            .I(N__16251));
    Odrv4 I__3463 (
            .O(N__16267),
            .I(\Lab_UT.de_cr_6_0 ));
    Odrv4 I__3462 (
            .O(N__16264),
            .I(\Lab_UT.de_cr_6_0 ));
    Odrv12 I__3461 (
            .O(N__16261),
            .I(\Lab_UT.de_cr_6_0 ));
    LocalMux I__3460 (
            .O(N__16256),
            .I(\Lab_UT.de_cr_6_0 ));
    LocalMux I__3459 (
            .O(N__16251),
            .I(\Lab_UT.de_cr_6_0 ));
    CascadeMux I__3458 (
            .O(N__16240),
            .I(\Lab_UT.g0_i_a5_1_3_cascade_ ));
    InMux I__3457 (
            .O(N__16237),
            .I(N__16234));
    LocalMux I__3456 (
            .O(N__16234),
            .I(\Lab_UT.scdp.a2b.N_9_1 ));
    CascadeMux I__3455 (
            .O(N__16231),
            .I(N__16227));
    CascadeMux I__3454 (
            .O(N__16230),
            .I(N__16224));
    InMux I__3453 (
            .O(N__16227),
            .I(N__16221));
    InMux I__3452 (
            .O(N__16224),
            .I(N__16218));
    LocalMux I__3451 (
            .O(N__16221),
            .I(\Lab_UT.scdp.a2b.g1_1_0_1 ));
    LocalMux I__3450 (
            .O(N__16218),
            .I(\Lab_UT.scdp.a2b.g1_1_0_1 ));
    InMux I__3449 (
            .O(N__16213),
            .I(N__16210));
    LocalMux I__3448 (
            .O(N__16210),
            .I(\Lab_UT.scctrl.g0_1_3_1 ));
    InMux I__3447 (
            .O(N__16207),
            .I(N__16204));
    LocalMux I__3446 (
            .O(N__16204),
            .I(N__16201));
    Span4Mux_v I__3445 (
            .O(N__16201),
            .I(N__16198));
    Span4Mux_s3_h I__3444 (
            .O(N__16198),
            .I(N__16195));
    Odrv4 I__3443 (
            .O(N__16195),
            .I(Lab_UT_dk_de_cr_12_1));
    CascadeMux I__3442 (
            .O(N__16192),
            .I(N__16189));
    InMux I__3441 (
            .O(N__16189),
            .I(N__16186));
    LocalMux I__3440 (
            .O(N__16186),
            .I(N__16181));
    InMux I__3439 (
            .O(N__16185),
            .I(N__16176));
    InMux I__3438 (
            .O(N__16184),
            .I(N__16176));
    Odrv12 I__3437 (
            .O(N__16181),
            .I(\ufifo.emptyB_0 ));
    LocalMux I__3436 (
            .O(N__16176),
            .I(\ufifo.emptyB_0 ));
    CascadeMux I__3435 (
            .O(N__16171),
            .I(N__16159));
    InMux I__3434 (
            .O(N__16170),
            .I(N__16156));
    InMux I__3433 (
            .O(N__16169),
            .I(N__16150));
    InMux I__3432 (
            .O(N__16168),
            .I(N__16150));
    InMux I__3431 (
            .O(N__16167),
            .I(N__16147));
    InMux I__3430 (
            .O(N__16166),
            .I(N__16143));
    InMux I__3429 (
            .O(N__16165),
            .I(N__16137));
    InMux I__3428 (
            .O(N__16164),
            .I(N__16137));
    InMux I__3427 (
            .O(N__16163),
            .I(N__16133));
    InMux I__3426 (
            .O(N__16162),
            .I(N__16128));
    InMux I__3425 (
            .O(N__16159),
            .I(N__16128));
    LocalMux I__3424 (
            .O(N__16156),
            .I(N__16125));
    InMux I__3423 (
            .O(N__16155),
            .I(N__16122));
    LocalMux I__3422 (
            .O(N__16150),
            .I(N__16119));
    LocalMux I__3421 (
            .O(N__16147),
            .I(N__16116));
    InMux I__3420 (
            .O(N__16146),
            .I(N__16113));
    LocalMux I__3419 (
            .O(N__16143),
            .I(N__16110));
    InMux I__3418 (
            .O(N__16142),
            .I(N__16107));
    LocalMux I__3417 (
            .O(N__16137),
            .I(N__16104));
    InMux I__3416 (
            .O(N__16136),
            .I(N__16101));
    LocalMux I__3415 (
            .O(N__16133),
            .I(N__16096));
    LocalMux I__3414 (
            .O(N__16128),
            .I(N__16096));
    Span4Mux_h I__3413 (
            .O(N__16125),
            .I(N__16089));
    LocalMux I__3412 (
            .O(N__16122),
            .I(N__16089));
    Span4Mux_h I__3411 (
            .O(N__16119),
            .I(N__16089));
    Span4Mux_h I__3410 (
            .O(N__16116),
            .I(N__16076));
    LocalMux I__3409 (
            .O(N__16113),
            .I(N__16076));
    Span4Mux_h I__3408 (
            .O(N__16110),
            .I(N__16076));
    LocalMux I__3407 (
            .O(N__16107),
            .I(N__16076));
    Span4Mux_h I__3406 (
            .O(N__16104),
            .I(N__16076));
    LocalMux I__3405 (
            .O(N__16101),
            .I(N__16076));
    Odrv4 I__3404 (
            .O(N__16096),
            .I(bu_rx_data_0));
    Odrv4 I__3403 (
            .O(N__16089),
            .I(bu_rx_data_0));
    Odrv4 I__3402 (
            .O(N__16076),
            .I(bu_rx_data_0));
    InMux I__3401 (
            .O(N__16069),
            .I(N__16066));
    LocalMux I__3400 (
            .O(N__16066),
            .I(N__16063));
    Odrv12 I__3399 (
            .O(N__16063),
            .I(\ufifo.tx_fsm.N_60_0 ));
    InMux I__3398 (
            .O(N__16060),
            .I(N__16057));
    LocalMux I__3397 (
            .O(N__16057),
            .I(N__16054));
    Span4Mux_h I__3396 (
            .O(N__16054),
            .I(N__16051));
    Odrv4 I__3395 (
            .O(N__16051),
            .I(\Lab_UT.scctrl.N_127_i_i_a6_0_0 ));
    InMux I__3394 (
            .O(N__16048),
            .I(N__16045));
    LocalMux I__3393 (
            .O(N__16045),
            .I(\Lab_UT.scctrl.N_11 ));
    InMux I__3392 (
            .O(N__16042),
            .I(N__16039));
    LocalMux I__3391 (
            .O(N__16039),
            .I(\Lab_UT.scctrl.G_21_i_a7_1_1 ));
    CascadeMux I__3390 (
            .O(N__16036),
            .I(N__16033));
    InMux I__3389 (
            .O(N__16033),
            .I(N__16030));
    LocalMux I__3388 (
            .O(N__16030),
            .I(N__16027));
    Odrv12 I__3387 (
            .O(N__16027),
            .I(\Lab_UT.m61_i_a2_2 ));
    InMux I__3386 (
            .O(N__16024),
            .I(N__16021));
    LocalMux I__3385 (
            .O(N__16021),
            .I(\Lab_UT.scctrl.g0_0_i_0_0 ));
    CascadeMux I__3384 (
            .O(N__16018),
            .I(\Lab_UT.N_5_cascade_ ));
    InMux I__3383 (
            .O(N__16015),
            .I(N__16012));
    LocalMux I__3382 (
            .O(N__16012),
            .I(\Lab_UT.g0_i_5 ));
    InMux I__3381 (
            .O(N__16009),
            .I(N__16006));
    LocalMux I__3380 (
            .O(N__16006),
            .I(\Lab_UT.scctrl.g0_14_mb_sn ));
    InMux I__3379 (
            .O(N__16003),
            .I(N__16000));
    LocalMux I__3378 (
            .O(N__16000),
            .I(G_23_0_0));
    CascadeMux I__3377 (
            .O(N__15997),
            .I(N__15994));
    InMux I__3376 (
            .O(N__15994),
            .I(N__15991));
    LocalMux I__3375 (
            .O(N__15991),
            .I(N__15988));
    Odrv4 I__3374 (
            .O(N__15988),
            .I(\Lab_UT.scctrl.N_12_1 ));
    InMux I__3373 (
            .O(N__15985),
            .I(N__15981));
    InMux I__3372 (
            .O(N__15984),
            .I(N__15978));
    LocalMux I__3371 (
            .O(N__15981),
            .I(\Lab_UT.scctrl.N_5_0 ));
    LocalMux I__3370 (
            .O(N__15978),
            .I(\Lab_UT.scctrl.N_5_0 ));
    InMux I__3369 (
            .O(N__15973),
            .I(N__15970));
    LocalMux I__3368 (
            .O(N__15970),
            .I(N__15967));
    Odrv4 I__3367 (
            .O(N__15967),
            .I(\Lab_UT.scctrl.g0_0_i_a8_3_1_0 ));
    CascadeMux I__3366 (
            .O(N__15964),
            .I(\Lab_UT.scctrl.g0_0_i_a8_2_1_0_cascade_ ));
    CascadeMux I__3365 (
            .O(N__15961),
            .I(\Lab_UT.scctrl.g0_0_i_3_0_cascade_ ));
    InMux I__3364 (
            .O(N__15958),
            .I(N__15955));
    LocalMux I__3363 (
            .O(N__15955),
            .I(\Lab_UT.scctrl.N_13 ));
    InMux I__3362 (
            .O(N__15952),
            .I(N__15949));
    LocalMux I__3361 (
            .O(N__15949),
            .I(\Lab_UT.scctrl.g0_i_1 ));
    InMux I__3360 (
            .O(N__15946),
            .I(N__15936));
    InMux I__3359 (
            .O(N__15945),
            .I(N__15936));
    InMux I__3358 (
            .O(N__15944),
            .I(N__15936));
    InMux I__3357 (
            .O(N__15943),
            .I(N__15933));
    LocalMux I__3356 (
            .O(N__15936),
            .I(\Lab_UT.scctrl.g0_0_i_2 ));
    LocalMux I__3355 (
            .O(N__15933),
            .I(\Lab_UT.scctrl.g0_0_i_2 ));
    CascadeMux I__3354 (
            .O(N__15928),
            .I(N__15925));
    InMux I__3353 (
            .O(N__15925),
            .I(N__15915));
    InMux I__3352 (
            .O(N__15924),
            .I(N__15915));
    InMux I__3351 (
            .O(N__15923),
            .I(N__15915));
    InMux I__3350 (
            .O(N__15922),
            .I(N__15911));
    LocalMux I__3349 (
            .O(N__15915),
            .I(N__15908));
    InMux I__3348 (
            .O(N__15914),
            .I(N__15905));
    LocalMux I__3347 (
            .O(N__15911),
            .I(\Lab_UT.scctrl.g0_16_mb_sn ));
    Odrv4 I__3346 (
            .O(N__15908),
            .I(\Lab_UT.scctrl.g0_16_mb_sn ));
    LocalMux I__3345 (
            .O(N__15905),
            .I(\Lab_UT.scctrl.g0_16_mb_sn ));
    CascadeMux I__3344 (
            .O(N__15898),
            .I(N__15892));
    CascadeMux I__3343 (
            .O(N__15897),
            .I(N__15888));
    InMux I__3342 (
            .O(N__15896),
            .I(N__15885));
    InMux I__3341 (
            .O(N__15895),
            .I(N__15878));
    InMux I__3340 (
            .O(N__15892),
            .I(N__15878));
    InMux I__3339 (
            .O(N__15891),
            .I(N__15878));
    InMux I__3338 (
            .O(N__15888),
            .I(N__15875));
    LocalMux I__3337 (
            .O(N__15885),
            .I(N__15868));
    LocalMux I__3336 (
            .O(N__15878),
            .I(N__15868));
    LocalMux I__3335 (
            .O(N__15875),
            .I(N__15868));
    Span4Mux_v I__3334 (
            .O(N__15868),
            .I(N__15865));
    Span4Mux_s3_h I__3333 (
            .O(N__15865),
            .I(N__15862));
    Odrv4 I__3332 (
            .O(N__15862),
            .I(\Lab_UT.scctrl.g0_16_mb_rn_0 ));
    InMux I__3331 (
            .O(N__15859),
            .I(N__15853));
    InMux I__3330 (
            .O(N__15858),
            .I(N__15848));
    InMux I__3329 (
            .O(N__15857),
            .I(N__15848));
    InMux I__3328 (
            .O(N__15856),
            .I(N__15845));
    LocalMux I__3327 (
            .O(N__15853),
            .I(\Lab_UT.scctrl.g0_0_i_3_0 ));
    LocalMux I__3326 (
            .O(N__15848),
            .I(\Lab_UT.scctrl.g0_0_i_3_0 ));
    LocalMux I__3325 (
            .O(N__15845),
            .I(\Lab_UT.scctrl.g0_0_i_3_0 ));
    InMux I__3324 (
            .O(N__15838),
            .I(N__15835));
    LocalMux I__3323 (
            .O(N__15835),
            .I(N__15831));
    InMux I__3322 (
            .O(N__15834),
            .I(N__15828));
    Span4Mux_h I__3321 (
            .O(N__15831),
            .I(N__15825));
    LocalMux I__3320 (
            .O(N__15828),
            .I(\Lab_UT.scdp.key0_5 ));
    Odrv4 I__3319 (
            .O(N__15825),
            .I(\Lab_UT.scdp.key0_5 ));
    InMux I__3318 (
            .O(N__15820),
            .I(N__15813));
    InMux I__3317 (
            .O(N__15819),
            .I(N__15813));
    InMux I__3316 (
            .O(N__15818),
            .I(N__15810));
    LocalMux I__3315 (
            .O(N__15813),
            .I(N__15806));
    LocalMux I__3314 (
            .O(N__15810),
            .I(N__15803));
    InMux I__3313 (
            .O(N__15809),
            .I(N__15800));
    Span4Mux_h I__3312 (
            .O(N__15806),
            .I(N__15793));
    Span4Mux_h I__3311 (
            .O(N__15803),
            .I(N__15793));
    LocalMux I__3310 (
            .O(N__15800),
            .I(N__15793));
    Odrv4 I__3309 (
            .O(N__15793),
            .I(\Lab_UT.scdp.a2b.N_53 ));
    CascadeMux I__3308 (
            .O(N__15790),
            .I(N__15786));
    CascadeMux I__3307 (
            .O(N__15789),
            .I(N__15783));
    InMux I__3306 (
            .O(N__15786),
            .I(N__15777));
    InMux I__3305 (
            .O(N__15783),
            .I(N__15777));
    InMux I__3304 (
            .O(N__15782),
            .I(N__15773));
    LocalMux I__3303 (
            .O(N__15777),
            .I(N__15768));
    InMux I__3302 (
            .O(N__15776),
            .I(N__15765));
    LocalMux I__3301 (
            .O(N__15773),
            .I(N__15762));
    InMux I__3300 (
            .O(N__15772),
            .I(N__15759));
    InMux I__3299 (
            .O(N__15771),
            .I(N__15755));
    Span4Mux_h I__3298 (
            .O(N__15768),
            .I(N__15747));
    LocalMux I__3297 (
            .O(N__15765),
            .I(N__15747));
    Span4Mux_v I__3296 (
            .O(N__15762),
            .I(N__15742));
    LocalMux I__3295 (
            .O(N__15759),
            .I(N__15742));
    InMux I__3294 (
            .O(N__15758),
            .I(N__15739));
    LocalMux I__3293 (
            .O(N__15755),
            .I(N__15736));
    InMux I__3292 (
            .O(N__15754),
            .I(N__15733));
    InMux I__3291 (
            .O(N__15753),
            .I(N__15728));
    InMux I__3290 (
            .O(N__15752),
            .I(N__15728));
    Span4Mux_v I__3289 (
            .O(N__15747),
            .I(N__15723));
    Span4Mux_h I__3288 (
            .O(N__15742),
            .I(N__15723));
    LocalMux I__3287 (
            .O(N__15739),
            .I(N__15720));
    Span4Mux_v I__3286 (
            .O(N__15736),
            .I(N__15717));
    LocalMux I__3285 (
            .O(N__15733),
            .I(bu_rx_data_1));
    LocalMux I__3284 (
            .O(N__15728),
            .I(bu_rx_data_1));
    Odrv4 I__3283 (
            .O(N__15723),
            .I(bu_rx_data_1));
    Odrv12 I__3282 (
            .O(N__15720),
            .I(bu_rx_data_1));
    Odrv4 I__3281 (
            .O(N__15717),
            .I(bu_rx_data_1));
    InMux I__3280 (
            .O(N__15706),
            .I(N__15697));
    InMux I__3279 (
            .O(N__15705),
            .I(N__15697));
    CascadeMux I__3278 (
            .O(N__15704),
            .I(N__15691));
    CascadeMux I__3277 (
            .O(N__15703),
            .I(N__15688));
    CascadeMux I__3276 (
            .O(N__15702),
            .I(N__15683));
    LocalMux I__3275 (
            .O(N__15697),
            .I(N__15677));
    InMux I__3274 (
            .O(N__15696),
            .I(N__15674));
    InMux I__3273 (
            .O(N__15695),
            .I(N__15671));
    InMux I__3272 (
            .O(N__15694),
            .I(N__15666));
    InMux I__3271 (
            .O(N__15691),
            .I(N__15666));
    InMux I__3270 (
            .O(N__15688),
            .I(N__15662));
    InMux I__3269 (
            .O(N__15687),
            .I(N__15659));
    InMux I__3268 (
            .O(N__15686),
            .I(N__15656));
    InMux I__3267 (
            .O(N__15683),
            .I(N__15653));
    InMux I__3266 (
            .O(N__15682),
            .I(N__15647));
    InMux I__3265 (
            .O(N__15681),
            .I(N__15642));
    InMux I__3264 (
            .O(N__15680),
            .I(N__15642));
    Span4Mux_v I__3263 (
            .O(N__15677),
            .I(N__15639));
    LocalMux I__3262 (
            .O(N__15674),
            .I(N__15636));
    LocalMux I__3261 (
            .O(N__15671),
            .I(N__15633));
    LocalMux I__3260 (
            .O(N__15666),
            .I(N__15630));
    InMux I__3259 (
            .O(N__15665),
            .I(N__15627));
    LocalMux I__3258 (
            .O(N__15662),
            .I(N__15624));
    LocalMux I__3257 (
            .O(N__15659),
            .I(N__15621));
    LocalMux I__3256 (
            .O(N__15656),
            .I(N__15618));
    LocalMux I__3255 (
            .O(N__15653),
            .I(N__15615));
    InMux I__3254 (
            .O(N__15652),
            .I(N__15612));
    InMux I__3253 (
            .O(N__15651),
            .I(N__15607));
    InMux I__3252 (
            .O(N__15650),
            .I(N__15607));
    LocalMux I__3251 (
            .O(N__15647),
            .I(N__15602));
    LocalMux I__3250 (
            .O(N__15642),
            .I(N__15602));
    Span4Mux_v I__3249 (
            .O(N__15639),
            .I(N__15593));
    Span4Mux_v I__3248 (
            .O(N__15636),
            .I(N__15593));
    Span4Mux_v I__3247 (
            .O(N__15633),
            .I(N__15593));
    Span4Mux_v I__3246 (
            .O(N__15630),
            .I(N__15593));
    LocalMux I__3245 (
            .O(N__15627),
            .I(N__15588));
    Span4Mux_h I__3244 (
            .O(N__15624),
            .I(N__15588));
    Span4Mux_v I__3243 (
            .O(N__15621),
            .I(N__15581));
    Span4Mux_v I__3242 (
            .O(N__15618),
            .I(N__15581));
    Span4Mux_s2_h I__3241 (
            .O(N__15615),
            .I(N__15581));
    LocalMux I__3240 (
            .O(N__15612),
            .I(bu_rx_data_2));
    LocalMux I__3239 (
            .O(N__15607),
            .I(bu_rx_data_2));
    Odrv12 I__3238 (
            .O(N__15602),
            .I(bu_rx_data_2));
    Odrv4 I__3237 (
            .O(N__15593),
            .I(bu_rx_data_2));
    Odrv4 I__3236 (
            .O(N__15588),
            .I(bu_rx_data_2));
    Odrv4 I__3235 (
            .O(N__15581),
            .I(bu_rx_data_2));
    InMux I__3234 (
            .O(N__15568),
            .I(N__15562));
    InMux I__3233 (
            .O(N__15567),
            .I(N__15562));
    LocalMux I__3232 (
            .O(N__15562),
            .I(N__15553));
    InMux I__3231 (
            .O(N__15561),
            .I(N__15550));
    InMux I__3230 (
            .O(N__15560),
            .I(N__15541));
    InMux I__3229 (
            .O(N__15559),
            .I(N__15541));
    InMux I__3228 (
            .O(N__15558),
            .I(N__15541));
    InMux I__3227 (
            .O(N__15557),
            .I(N__15541));
    InMux I__3226 (
            .O(N__15556),
            .I(N__15538));
    Odrv4 I__3225 (
            .O(N__15553),
            .I(\Lab_UT.scdp.binValD_2 ));
    LocalMux I__3224 (
            .O(N__15550),
            .I(\Lab_UT.scdp.binValD_2 ));
    LocalMux I__3223 (
            .O(N__15541),
            .I(\Lab_UT.scdp.binValD_2 ));
    LocalMux I__3222 (
            .O(N__15538),
            .I(\Lab_UT.scdp.binValD_2 ));
    InMux I__3221 (
            .O(N__15529),
            .I(N__15525));
    InMux I__3220 (
            .O(N__15528),
            .I(N__15522));
    LocalMux I__3219 (
            .O(N__15525),
            .I(N__15519));
    LocalMux I__3218 (
            .O(N__15522),
            .I(N__15514));
    Span4Mux_v I__3217 (
            .O(N__15519),
            .I(N__15514));
    Odrv4 I__3216 (
            .O(N__15514),
            .I(\Lab_UT.scdp.key0_6 ));
    InMux I__3215 (
            .O(N__15511),
            .I(N__15506));
    InMux I__3214 (
            .O(N__15510),
            .I(N__15503));
    CascadeMux I__3213 (
            .O(N__15509),
            .I(N__15500));
    LocalMux I__3212 (
            .O(N__15506),
            .I(N__15494));
    LocalMux I__3211 (
            .O(N__15503),
            .I(N__15491));
    InMux I__3210 (
            .O(N__15500),
            .I(N__15482));
    InMux I__3209 (
            .O(N__15499),
            .I(N__15482));
    InMux I__3208 (
            .O(N__15498),
            .I(N__15482));
    InMux I__3207 (
            .O(N__15497),
            .I(N__15479));
    Span4Mux_v I__3206 (
            .O(N__15494),
            .I(N__15474));
    Span4Mux_v I__3205 (
            .O(N__15491),
            .I(N__15474));
    InMux I__3204 (
            .O(N__15490),
            .I(N__15469));
    InMux I__3203 (
            .O(N__15489),
            .I(N__15469));
    LocalMux I__3202 (
            .O(N__15482),
            .I(N__15464));
    LocalMux I__3201 (
            .O(N__15479),
            .I(N__15464));
    Span4Mux_s3_h I__3200 (
            .O(N__15474),
            .I(N__15461));
    LocalMux I__3199 (
            .O(N__15469),
            .I(\Lab_UT.scdp.binValD_0 ));
    Odrv12 I__3198 (
            .O(N__15464),
            .I(\Lab_UT.scdp.binValD_0 ));
    Odrv4 I__3197 (
            .O(N__15461),
            .I(\Lab_UT.scdp.binValD_0 ));
    InMux I__3196 (
            .O(N__15454),
            .I(N__15451));
    LocalMux I__3195 (
            .O(N__15451),
            .I(N__15448));
    Span4Mux_v I__3194 (
            .O(N__15448),
            .I(N__15444));
    InMux I__3193 (
            .O(N__15447),
            .I(N__15441));
    Span4Mux_s2_v I__3192 (
            .O(N__15444),
            .I(N__15438));
    LocalMux I__3191 (
            .O(N__15441),
            .I(\Lab_UT.scdp.key0_4 ));
    Odrv4 I__3190 (
            .O(N__15438),
            .I(\Lab_UT.scdp.key0_4 ));
    InMux I__3189 (
            .O(N__15433),
            .I(N__15426));
    InMux I__3188 (
            .O(N__15432),
            .I(N__15417));
    InMux I__3187 (
            .O(N__15431),
            .I(N__15417));
    InMux I__3186 (
            .O(N__15430),
            .I(N__15417));
    InMux I__3185 (
            .O(N__15429),
            .I(N__15417));
    LocalMux I__3184 (
            .O(N__15426),
            .I(\Lab_UT.state_ret_RNIUV0941_0 ));
    LocalMux I__3183 (
            .O(N__15417),
            .I(\Lab_UT.state_ret_RNIUV0941_0 ));
    InMux I__3182 (
            .O(N__15412),
            .I(N__15408));
    CascadeMux I__3181 (
            .O(N__15411),
            .I(N__15405));
    LocalMux I__3180 (
            .O(N__15408),
            .I(N__15402));
    InMux I__3179 (
            .O(N__15405),
            .I(N__15399));
    Span4Mux_h I__3178 (
            .O(N__15402),
            .I(N__15396));
    LocalMux I__3177 (
            .O(N__15399),
            .I(\Lab_UT.scdp.key0_7 ));
    Odrv4 I__3176 (
            .O(N__15396),
            .I(\Lab_UT.scdp.key0_7 ));
    CascadeMux I__3175 (
            .O(N__15391),
            .I(N__15387));
    CascadeMux I__3174 (
            .O(N__15390),
            .I(N__15380));
    InMux I__3173 (
            .O(N__15387),
            .I(N__15369));
    InMux I__3172 (
            .O(N__15386),
            .I(N__15369));
    InMux I__3171 (
            .O(N__15385),
            .I(N__15369));
    InMux I__3170 (
            .O(N__15384),
            .I(N__15369));
    InMux I__3169 (
            .O(N__15383),
            .I(N__15369));
    InMux I__3168 (
            .O(N__15380),
            .I(N__15366));
    LocalMux I__3167 (
            .O(N__15369),
            .I(N__15361));
    LocalMux I__3166 (
            .O(N__15366),
            .I(N__15358));
    InMux I__3165 (
            .O(N__15365),
            .I(N__15353));
    InMux I__3164 (
            .O(N__15364),
            .I(N__15353));
    Span4Mux_s2_v I__3163 (
            .O(N__15361),
            .I(N__15350));
    Odrv12 I__3162 (
            .O(N__15358),
            .I(\Lab_UT.scdp.binValD_1 ));
    LocalMux I__3161 (
            .O(N__15353),
            .I(\Lab_UT.scdp.binValD_1 ));
    Odrv4 I__3160 (
            .O(N__15350),
            .I(\Lab_UT.scdp.binValD_1 ));
    InMux I__3159 (
            .O(N__15343),
            .I(N__15340));
    LocalMux I__3158 (
            .O(N__15340),
            .I(N__15336));
    InMux I__3157 (
            .O(N__15339),
            .I(N__15333));
    Span4Mux_h I__3156 (
            .O(N__15336),
            .I(N__15330));
    LocalMux I__3155 (
            .O(N__15333),
            .I(\Lab_UT.scdp.key0_1 ));
    Odrv4 I__3154 (
            .O(N__15330),
            .I(\Lab_UT.scdp.key0_1 ));
    InMux I__3153 (
            .O(N__15325),
            .I(N__15318));
    InMux I__3152 (
            .O(N__15324),
            .I(N__15313));
    InMux I__3151 (
            .O(N__15323),
            .I(N__15306));
    InMux I__3150 (
            .O(N__15322),
            .I(N__15306));
    InMux I__3149 (
            .O(N__15321),
            .I(N__15306));
    LocalMux I__3148 (
            .O(N__15318),
            .I(N__15303));
    InMux I__3147 (
            .O(N__15317),
            .I(N__15298));
    InMux I__3146 (
            .O(N__15316),
            .I(N__15298));
    LocalMux I__3145 (
            .O(N__15313),
            .I(N__15291));
    LocalMux I__3144 (
            .O(N__15306),
            .I(N__15291));
    Span4Mux_s2_v I__3143 (
            .O(N__15303),
            .I(N__15291));
    LocalMux I__3142 (
            .O(N__15298),
            .I(\Lab_UT.scdp.binValD_3 ));
    Odrv4 I__3141 (
            .O(N__15291),
            .I(\Lab_UT.scdp.binValD_3 ));
    CascadeMux I__3140 (
            .O(N__15286),
            .I(N__15283));
    InMux I__3139 (
            .O(N__15283),
            .I(N__15269));
    CascadeMux I__3138 (
            .O(N__15282),
            .I(N__15266));
    CascadeMux I__3137 (
            .O(N__15281),
            .I(N__15262));
    CascadeMux I__3136 (
            .O(N__15280),
            .I(N__15259));
    CascadeMux I__3135 (
            .O(N__15279),
            .I(N__15256));
    CascadeMux I__3134 (
            .O(N__15278),
            .I(N__15253));
    CascadeMux I__3133 (
            .O(N__15277),
            .I(N__15244));
    CascadeMux I__3132 (
            .O(N__15276),
            .I(N__15241));
    CascadeMux I__3131 (
            .O(N__15275),
            .I(N__15237));
    CascadeMux I__3130 (
            .O(N__15274),
            .I(N__15234));
    CascadeMux I__3129 (
            .O(N__15273),
            .I(N__15225));
    CascadeMux I__3128 (
            .O(N__15272),
            .I(N__15220));
    LocalMux I__3127 (
            .O(N__15269),
            .I(N__15217));
    InMux I__3126 (
            .O(N__15266),
            .I(N__15214));
    InMux I__3125 (
            .O(N__15265),
            .I(N__15203));
    InMux I__3124 (
            .O(N__15262),
            .I(N__15203));
    InMux I__3123 (
            .O(N__15259),
            .I(N__15203));
    InMux I__3122 (
            .O(N__15256),
            .I(N__15203));
    InMux I__3121 (
            .O(N__15253),
            .I(N__15203));
    CascadeMux I__3120 (
            .O(N__15252),
            .I(N__15200));
    CascadeMux I__3119 (
            .O(N__15251),
            .I(N__15197));
    CascadeMux I__3118 (
            .O(N__15250),
            .I(N__15194));
    CascadeMux I__3117 (
            .O(N__15249),
            .I(N__15191));
    CascadeMux I__3116 (
            .O(N__15248),
            .I(N__15188));
    CascadeMux I__3115 (
            .O(N__15247),
            .I(N__15185));
    InMux I__3114 (
            .O(N__15244),
            .I(N__15175));
    InMux I__3113 (
            .O(N__15241),
            .I(N__15175));
    InMux I__3112 (
            .O(N__15240),
            .I(N__15175));
    InMux I__3111 (
            .O(N__15237),
            .I(N__15158));
    InMux I__3110 (
            .O(N__15234),
            .I(N__15158));
    InMux I__3109 (
            .O(N__15233),
            .I(N__15158));
    InMux I__3108 (
            .O(N__15232),
            .I(N__15158));
    InMux I__3107 (
            .O(N__15231),
            .I(N__15158));
    InMux I__3106 (
            .O(N__15230),
            .I(N__15158));
    InMux I__3105 (
            .O(N__15229),
            .I(N__15158));
    InMux I__3104 (
            .O(N__15228),
            .I(N__15158));
    InMux I__3103 (
            .O(N__15225),
            .I(N__15151));
    InMux I__3102 (
            .O(N__15224),
            .I(N__15151));
    InMux I__3101 (
            .O(N__15223),
            .I(N__15151));
    InMux I__3100 (
            .O(N__15220),
            .I(N__15148));
    Span4Mux_v I__3099 (
            .O(N__15217),
            .I(N__15143));
    LocalMux I__3098 (
            .O(N__15214),
            .I(N__15143));
    LocalMux I__3097 (
            .O(N__15203),
            .I(N__15140));
    InMux I__3096 (
            .O(N__15200),
            .I(N__15135));
    InMux I__3095 (
            .O(N__15197),
            .I(N__15135));
    InMux I__3094 (
            .O(N__15194),
            .I(N__15132));
    InMux I__3093 (
            .O(N__15191),
            .I(N__15129));
    InMux I__3092 (
            .O(N__15188),
            .I(N__15118));
    InMux I__3091 (
            .O(N__15185),
            .I(N__15118));
    InMux I__3090 (
            .O(N__15184),
            .I(N__15118));
    InMux I__3089 (
            .O(N__15183),
            .I(N__15118));
    InMux I__3088 (
            .O(N__15182),
            .I(N__15118));
    LocalMux I__3087 (
            .O(N__15175),
            .I(N__15115));
    LocalMux I__3086 (
            .O(N__15158),
            .I(N__15112));
    LocalMux I__3085 (
            .O(N__15151),
            .I(N__15109));
    LocalMux I__3084 (
            .O(N__15148),
            .I(N__15104));
    Span4Mux_h I__3083 (
            .O(N__15143),
            .I(N__15104));
    Span4Mux_h I__3082 (
            .O(N__15140),
            .I(N__15101));
    LocalMux I__3081 (
            .O(N__15135),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    LocalMux I__3080 (
            .O(N__15132),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    LocalMux I__3079 (
            .O(N__15129),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    LocalMux I__3078 (
            .O(N__15118),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    Odrv4 I__3077 (
            .O(N__15115),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    Odrv12 I__3076 (
            .O(N__15112),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    Odrv12 I__3075 (
            .O(N__15109),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    Odrv4 I__3074 (
            .O(N__15104),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    Odrv4 I__3073 (
            .O(N__15101),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    InMux I__3072 (
            .O(N__15082),
            .I(N__15078));
    InMux I__3071 (
            .O(N__15081),
            .I(N__15072));
    LocalMux I__3070 (
            .O(N__15078),
            .I(N__15069));
    InMux I__3069 (
            .O(N__15077),
            .I(N__15066));
    InMux I__3068 (
            .O(N__15076),
            .I(N__15061));
    InMux I__3067 (
            .O(N__15075),
            .I(N__15061));
    LocalMux I__3066 (
            .O(N__15072),
            .I(\Lab_UT.state_0_RNIKFK051_0_1 ));
    Odrv4 I__3065 (
            .O(N__15069),
            .I(\Lab_UT.state_0_RNIKFK051_0_1 ));
    LocalMux I__3064 (
            .O(N__15066),
            .I(\Lab_UT.state_0_RNIKFK051_0_1 ));
    LocalMux I__3063 (
            .O(N__15061),
            .I(\Lab_UT.state_0_RNIKFK051_0_1 ));
    InMux I__3062 (
            .O(N__15052),
            .I(N__15049));
    LocalMux I__3061 (
            .O(N__15049),
            .I(N__15045));
    InMux I__3060 (
            .O(N__15048),
            .I(N__15042));
    Span4Mux_h I__3059 (
            .O(N__15045),
            .I(N__15039));
    LocalMux I__3058 (
            .O(N__15042),
            .I(\Lab_UT.scdp.key0_3 ));
    Odrv4 I__3057 (
            .O(N__15039),
            .I(\Lab_UT.scdp.key0_3 ));
    InMux I__3056 (
            .O(N__15034),
            .I(N__15031));
    LocalMux I__3055 (
            .O(N__15031),
            .I(N__15027));
    InMux I__3054 (
            .O(N__15030),
            .I(N__15024));
    Span4Mux_v I__3053 (
            .O(N__15027),
            .I(N__15021));
    LocalMux I__3052 (
            .O(N__15024),
            .I(N__15018));
    Odrv4 I__3051 (
            .O(N__15021),
            .I(\Lab_UT.scctrl.next_state74 ));
    Odrv4 I__3050 (
            .O(N__15018),
            .I(\Lab_UT.scctrl.next_state74 ));
    CascadeMux I__3049 (
            .O(N__15013),
            .I(N__15010));
    InMux I__3048 (
            .O(N__15010),
            .I(N__15007));
    LocalMux I__3047 (
            .O(N__15007),
            .I(N__15004));
    Odrv12 I__3046 (
            .O(N__15004),
            .I(\Lab_UT.scctrl.N_7_1 ));
    InMux I__3045 (
            .O(N__15001),
            .I(N__14998));
    LocalMux I__3044 (
            .O(N__14998),
            .I(\Lab_UT.scctrl.N_223_2 ));
    InMux I__3043 (
            .O(N__14995),
            .I(N__14992));
    LocalMux I__3042 (
            .O(N__14992),
            .I(\Lab_UT.scctrl.next_state73 ));
    CascadeMux I__3041 (
            .O(N__14989),
            .I(\Lab_UT.scctrl.next_state73_cascade_ ));
    InMux I__3040 (
            .O(N__14986),
            .I(N__14973));
    InMux I__3039 (
            .O(N__14985),
            .I(N__14973));
    InMux I__3038 (
            .O(N__14984),
            .I(N__14973));
    InMux I__3037 (
            .O(N__14983),
            .I(N__14970));
    InMux I__3036 (
            .O(N__14982),
            .I(N__14967));
    InMux I__3035 (
            .O(N__14981),
            .I(N__14964));
    InMux I__3034 (
            .O(N__14980),
            .I(N__14961));
    LocalMux I__3033 (
            .O(N__14973),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i ));
    LocalMux I__3032 (
            .O(N__14970),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i ));
    LocalMux I__3031 (
            .O(N__14967),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i ));
    LocalMux I__3030 (
            .O(N__14964),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i ));
    LocalMux I__3029 (
            .O(N__14961),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i ));
    CascadeMux I__3028 (
            .O(N__14950),
            .I(\Lab_UT.state_ret_3_RNII68F41_0_cascade_ ));
    InMux I__3027 (
            .O(N__14947),
            .I(N__14944));
    LocalMux I__3026 (
            .O(N__14944),
            .I(N__14940));
    InMux I__3025 (
            .O(N__14943),
            .I(N__14937));
    Span4Mux_h I__3024 (
            .O(N__14940),
            .I(N__14934));
    LocalMux I__3023 (
            .O(N__14937),
            .I(\Lab_UT.scdp.key2_0 ));
    Odrv4 I__3022 (
            .O(N__14934),
            .I(\Lab_UT.scdp.key2_0 ));
    InMux I__3021 (
            .O(N__14929),
            .I(N__14925));
    InMux I__3020 (
            .O(N__14928),
            .I(N__14922));
    LocalMux I__3019 (
            .O(N__14925),
            .I(N__14919));
    LocalMux I__3018 (
            .O(N__14922),
            .I(N__14914));
    Span4Mux_h I__3017 (
            .O(N__14919),
            .I(N__14914));
    Odrv4 I__3016 (
            .O(N__14914),
            .I(\Lab_UT.scdp.key2_1 ));
    InMux I__3015 (
            .O(N__14911),
            .I(N__14905));
    InMux I__3014 (
            .O(N__14910),
            .I(N__14898));
    InMux I__3013 (
            .O(N__14909),
            .I(N__14898));
    InMux I__3012 (
            .O(N__14908),
            .I(N__14898));
    LocalMux I__3011 (
            .O(N__14905),
            .I(\Lab_UT.state_ret_3_RNII68F41_0 ));
    LocalMux I__3010 (
            .O(N__14898),
            .I(\Lab_UT.state_ret_3_RNII68F41_0 ));
    InMux I__3009 (
            .O(N__14893),
            .I(N__14890));
    LocalMux I__3008 (
            .O(N__14890),
            .I(N__14887));
    Span4Mux_v I__3007 (
            .O(N__14887),
            .I(N__14883));
    InMux I__3006 (
            .O(N__14886),
            .I(N__14880));
    Span4Mux_h I__3005 (
            .O(N__14883),
            .I(N__14877));
    LocalMux I__3004 (
            .O(N__14880),
            .I(\Lab_UT.scdp.key2_2 ));
    Odrv4 I__3003 (
            .O(N__14877),
            .I(\Lab_UT.scdp.key2_2 ));
    InMux I__3002 (
            .O(N__14872),
            .I(N__14869));
    LocalMux I__3001 (
            .O(N__14869),
            .I(N__14863));
    InMux I__3000 (
            .O(N__14868),
            .I(N__14856));
    InMux I__2999 (
            .O(N__14867),
            .I(N__14856));
    InMux I__2998 (
            .O(N__14866),
            .I(N__14856));
    Span4Mux_v I__2997 (
            .O(N__14863),
            .I(N__14849));
    LocalMux I__2996 (
            .O(N__14856),
            .I(N__14849));
    InMux I__2995 (
            .O(N__14855),
            .I(N__14846));
    CascadeMux I__2994 (
            .O(N__14854),
            .I(N__14841));
    Span4Mux_h I__2993 (
            .O(N__14849),
            .I(N__14838));
    LocalMux I__2992 (
            .O(N__14846),
            .I(N__14835));
    InMux I__2991 (
            .O(N__14845),
            .I(N__14830));
    InMux I__2990 (
            .O(N__14844),
            .I(N__14830));
    InMux I__2989 (
            .O(N__14841),
            .I(N__14827));
    Odrv4 I__2988 (
            .O(N__14838),
            .I(bu_rx_data_i_3_1));
    Odrv4 I__2987 (
            .O(N__14835),
            .I(bu_rx_data_i_3_1));
    LocalMux I__2986 (
            .O(N__14830),
            .I(bu_rx_data_i_3_1));
    LocalMux I__2985 (
            .O(N__14827),
            .I(bu_rx_data_i_3_1));
    CascadeMux I__2984 (
            .O(N__14818),
            .I(N__14815));
    InMux I__2983 (
            .O(N__14815),
            .I(N__14809));
    InMux I__2982 (
            .O(N__14814),
            .I(N__14809));
    LocalMux I__2981 (
            .O(N__14809),
            .I(\Lab_UT.scctrl.g0_i_2_0 ));
    InMux I__2980 (
            .O(N__14806),
            .I(N__14802));
    InMux I__2979 (
            .O(N__14805),
            .I(N__14799));
    LocalMux I__2978 (
            .O(N__14802),
            .I(\Lab_UT.scctrl.next_state_rst_0_3_N_6_1 ));
    LocalMux I__2977 (
            .O(N__14799),
            .I(\Lab_UT.scctrl.next_state_rst_0_3_N_6_1 ));
    CEMux I__2976 (
            .O(N__14794),
            .I(N__14788));
    CEMux I__2975 (
            .O(N__14793),
            .I(N__14785));
    CEMux I__2974 (
            .O(N__14792),
            .I(N__14782));
    CEMux I__2973 (
            .O(N__14791),
            .I(N__14779));
    LocalMux I__2972 (
            .O(N__14788),
            .I(N__14776));
    LocalMux I__2971 (
            .O(N__14785),
            .I(N__14773));
    LocalMux I__2970 (
            .O(N__14782),
            .I(N__14770));
    LocalMux I__2969 (
            .O(N__14779),
            .I(N__14767));
    Span4Mux_v I__2968 (
            .O(N__14776),
            .I(N__14762));
    Span4Mux_h I__2967 (
            .O(N__14773),
            .I(N__14762));
    Span4Mux_v I__2966 (
            .O(N__14770),
            .I(N__14757));
    Span4Mux_v I__2965 (
            .O(N__14767),
            .I(N__14757));
    Odrv4 I__2964 (
            .O(N__14762),
            .I(\Lab_UT.g0_3_0 ));
    Odrv4 I__2963 (
            .O(N__14757),
            .I(\Lab_UT.g0_3_0 ));
    CascadeMux I__2962 (
            .O(N__14752),
            .I(N__14749));
    InMux I__2961 (
            .O(N__14749),
            .I(N__14746));
    LocalMux I__2960 (
            .O(N__14746),
            .I(\Lab_UT.scctrl.g0_i_a8_3_0 ));
    InMux I__2959 (
            .O(N__14743),
            .I(N__14740));
    LocalMux I__2958 (
            .O(N__14740),
            .I(\Lab_UT.scctrl.N_6_3 ));
    CascadeMux I__2957 (
            .O(N__14737),
            .I(\Lab_UT.scctrl.g0_i_1_1_cascade_ ));
    CascadeMux I__2956 (
            .O(N__14734),
            .I(\Lab_UT.scctrl.next_state_1_0_1_3_cascade_ ));
    InMux I__2955 (
            .O(N__14731),
            .I(N__14728));
    LocalMux I__2954 (
            .O(N__14728),
            .I(N__14724));
    InMux I__2953 (
            .O(N__14727),
            .I(N__14721));
    Odrv4 I__2952 (
            .O(N__14724),
            .I(\Lab_UT.scctrl.next_state75 ));
    LocalMux I__2951 (
            .O(N__14721),
            .I(\Lab_UT.scctrl.next_state75 ));
    CascadeMux I__2950 (
            .O(N__14716),
            .I(\Lab_UT.scctrl.next_state_rst_1_3_1_cascade_ ));
    InMux I__2949 (
            .O(N__14713),
            .I(N__14710));
    LocalMux I__2948 (
            .O(N__14710),
            .I(N__14707));
    Odrv4 I__2947 (
            .O(N__14707),
            .I(\Lab_UT.next_state_rst_1_3 ));
    CascadeMux I__2946 (
            .O(N__14704),
            .I(\Lab_UT.next_state_rst_1_3_cascade_ ));
    InMux I__2945 (
            .O(N__14701),
            .I(N__14697));
    InMux I__2944 (
            .O(N__14700),
            .I(N__14694));
    LocalMux I__2943 (
            .O(N__14697),
            .I(N__14691));
    LocalMux I__2942 (
            .O(N__14694),
            .I(N__14688));
    Span4Mux_h I__2941 (
            .O(N__14691),
            .I(N__14685));
    Odrv12 I__2940 (
            .O(N__14688),
            .I(\Lab_UT.scctrl.N_166_0 ));
    Odrv4 I__2939 (
            .O(N__14685),
            .I(\Lab_UT.scctrl.N_166_0 ));
    CascadeMux I__2938 (
            .O(N__14680),
            .I(\Lab_UT.scctrl.next_state_rst_1_cascade_ ));
    CascadeMux I__2937 (
            .O(N__14677),
            .I(N__14673));
    InMux I__2936 (
            .O(N__14676),
            .I(N__14669));
    InMux I__2935 (
            .O(N__14673),
            .I(N__14666));
    IoInMux I__2934 (
            .O(N__14672),
            .I(N__14663));
    LocalMux I__2933 (
            .O(N__14669),
            .I(N__14660));
    LocalMux I__2932 (
            .O(N__14666),
            .I(N__14657));
    LocalMux I__2931 (
            .O(N__14663),
            .I(N__14654));
    Span4Mux_v I__2930 (
            .O(N__14660),
            .I(N__14651));
    Span4Mux_h I__2929 (
            .O(N__14657),
            .I(N__14648));
    Odrv12 I__2928 (
            .O(N__14654),
            .I(led_c_2));
    Odrv4 I__2927 (
            .O(N__14651),
            .I(led_c_2));
    Odrv4 I__2926 (
            .O(N__14648),
            .I(led_c_2));
    InMux I__2925 (
            .O(N__14641),
            .I(N__14638));
    LocalMux I__2924 (
            .O(N__14638),
            .I(N__14635));
    Span4Mux_v I__2923 (
            .O(N__14635),
            .I(N__14632));
    Odrv4 I__2922 (
            .O(N__14632),
            .I(\Lab_UT.scctrl.g0_17_N_4LZ0Z5 ));
    CascadeMux I__2921 (
            .O(N__14629),
            .I(\Lab_UT.scctrl.next_state_rst_0_3_N_6_1_cascade_ ));
    CascadeMux I__2920 (
            .O(N__14626),
            .I(\Lab_UT.scctrl.g0_i_2_0_cascade_ ));
    InMux I__2919 (
            .O(N__14623),
            .I(N__14617));
    InMux I__2918 (
            .O(N__14622),
            .I(N__14617));
    LocalMux I__2917 (
            .O(N__14617),
            .I(\Lab_UT.scctrl.next_state_rst_0 ));
    CascadeMux I__2916 (
            .O(N__14614),
            .I(\Lab_UT.scctrl.g0_1_1_cascade_ ));
    InMux I__2915 (
            .O(N__14611),
            .I(N__14608));
    LocalMux I__2914 (
            .O(N__14608),
            .I(\Lab_UT.scctrl.g0_2_0 ));
    InMux I__2913 (
            .O(N__14605),
            .I(N__14602));
    LocalMux I__2912 (
            .O(N__14602),
            .I(N__14599));
    Odrv4 I__2911 (
            .O(N__14599),
            .I(\Lab_UT.scctrl.N_12_0 ));
    InMux I__2910 (
            .O(N__14596),
            .I(N__14593));
    LocalMux I__2909 (
            .O(N__14593),
            .I(\Lab_UT.scctrl.g0_i_1_0 ));
    CascadeMux I__2908 (
            .O(N__14590),
            .I(\Lab_UT.scctrl.g0_i_3_0_cascade_ ));
    InMux I__2907 (
            .O(N__14587),
            .I(N__14584));
    LocalMux I__2906 (
            .O(N__14584),
            .I(N__14581));
    Odrv4 I__2905 (
            .O(N__14581),
            .I(\Lab_UT.scctrl.un6_sccDecrypt_0 ));
    CascadeMux I__2904 (
            .O(N__14578),
            .I(\Lab_UT.scctrl.g1_1_0_cascade_ ));
    InMux I__2903 (
            .O(N__14575),
            .I(N__14572));
    LocalMux I__2902 (
            .O(N__14572),
            .I(\Lab_UT.scctrl.g2_0 ));
    CascadeMux I__2901 (
            .O(N__14569),
            .I(\Lab_UT.scctrl.g0_1_2_cascade_ ));
    InMux I__2900 (
            .O(N__14566),
            .I(N__14563));
    LocalMux I__2899 (
            .O(N__14563),
            .I(\Lab_UT.scctrl.g0_8_0 ));
    InMux I__2898 (
            .O(N__14560),
            .I(N__14557));
    LocalMux I__2897 (
            .O(N__14557),
            .I(\Lab_UT.scdp.a2b.g1_1_o2_0Z0Z_0 ));
    CascadeMux I__2896 (
            .O(N__14554),
            .I(\Lab_UT.scdp.a2b.N_6_1_cascade_ ));
    InMux I__2895 (
            .O(N__14551),
            .I(N__14548));
    LocalMux I__2894 (
            .O(N__14548),
            .I(\Lab_UT.scdp.a2b.g0_3_a3_0Z0Z_3 ));
    InMux I__2893 (
            .O(N__14545),
            .I(N__14542));
    LocalMux I__2892 (
            .O(N__14542),
            .I(N__14539));
    Span4Mux_h I__2891 (
            .O(N__14539),
            .I(N__14533));
    InMux I__2890 (
            .O(N__14538),
            .I(N__14526));
    InMux I__2889 (
            .O(N__14537),
            .I(N__14526));
    InMux I__2888 (
            .O(N__14536),
            .I(N__14526));
    Odrv4 I__2887 (
            .O(N__14533),
            .I(\Lab_UT.N_190 ));
    LocalMux I__2886 (
            .O(N__14526),
            .I(\Lab_UT.N_190 ));
    InMux I__2885 (
            .O(N__14521),
            .I(N__14518));
    LocalMux I__2884 (
            .O(N__14518),
            .I(N__14515));
    Span4Mux_h I__2883 (
            .O(N__14515),
            .I(N__14512));
    Odrv4 I__2882 (
            .O(N__14512),
            .I(\Lab_UT.scctrl.N_6_3_0 ));
    CascadeMux I__2881 (
            .O(N__14509),
            .I(N_127_i_i_1_cascade_));
    InMux I__2880 (
            .O(N__14506),
            .I(N__14503));
    LocalMux I__2879 (
            .O(N__14503),
            .I(N__14500));
    Odrv4 I__2878 (
            .O(N__14500),
            .I(\Lab_UT.scctrl.N_11_0 ));
    InMux I__2877 (
            .O(N__14497),
            .I(N__14494));
    LocalMux I__2876 (
            .O(N__14494),
            .I(\Lab_UT.N_166_0_0 ));
    InMux I__2875 (
            .O(N__14491),
            .I(N__14488));
    LocalMux I__2874 (
            .O(N__14488),
            .I(\Lab_UT.scctrl.N_127_i_i_3 ));
    CascadeMux I__2873 (
            .O(N__14485),
            .I(\Lab_UT.g1_i_a4_0_2_cascade_ ));
    CascadeMux I__2872 (
            .O(N__14482),
            .I(N__14479));
    InMux I__2871 (
            .O(N__14479),
            .I(N__14476));
    LocalMux I__2870 (
            .O(N__14476),
            .I(N__14470));
    InMux I__2869 (
            .O(N__14475),
            .I(N__14467));
    InMux I__2868 (
            .O(N__14474),
            .I(N__14464));
    InMux I__2867 (
            .O(N__14473),
            .I(N__14461));
    Span4Mux_v I__2866 (
            .O(N__14470),
            .I(N__14452));
    LocalMux I__2865 (
            .O(N__14467),
            .I(N__14452));
    LocalMux I__2864 (
            .O(N__14464),
            .I(N__14452));
    LocalMux I__2863 (
            .O(N__14461),
            .I(N__14452));
    Odrv4 I__2862 (
            .O(N__14452),
            .I(\Lab_UT.next_state_3 ));
    CascadeMux I__2861 (
            .O(N__14449),
            .I(\Lab_UT.g0_3_a3_0_4_cascade_ ));
    CascadeMux I__2860 (
            .O(N__14446),
            .I(\Lab_UT.scctrl.g0_0_i_2_cascade_ ));
    CascadeMux I__2859 (
            .O(N__14443),
            .I(N__14439));
    InMux I__2858 (
            .O(N__14442),
            .I(N__14434));
    InMux I__2857 (
            .O(N__14439),
            .I(N__14434));
    LocalMux I__2856 (
            .O(N__14434),
            .I(N__14430));
    InMux I__2855 (
            .O(N__14433),
            .I(N__14427));
    Span4Mux_h I__2854 (
            .O(N__14430),
            .I(N__14424));
    LocalMux I__2853 (
            .O(N__14427),
            .I(N__14421));
    Span4Mux_v I__2852 (
            .O(N__14424),
            .I(N__14418));
    Span4Mux_v I__2851 (
            .O(N__14421),
            .I(N__14415));
    Odrv4 I__2850 (
            .O(N__14418),
            .I(\Lab_UT.scctrl.state_i_3_fast_0 ));
    Odrv4 I__2849 (
            .O(N__14415),
            .I(\Lab_UT.scctrl.state_i_3_fast_0 ));
    InMux I__2848 (
            .O(N__14410),
            .I(N__14407));
    LocalMux I__2847 (
            .O(N__14407),
            .I(\Lab_UT.scctrl.g0_i_1_1_0 ));
    InMux I__2846 (
            .O(N__14404),
            .I(N__14401));
    LocalMux I__2845 (
            .O(N__14401),
            .I(N__14398));
    Span4Mux_h I__2844 (
            .O(N__14398),
            .I(N__14395));
    Odrv4 I__2843 (
            .O(N__14395),
            .I(\Lab_UT.scdp.a2b.N_6_0 ));
    InMux I__2842 (
            .O(N__14392),
            .I(N__14389));
    LocalMux I__2841 (
            .O(N__14389),
            .I(N__14386));
    Span4Mux_v I__2840 (
            .O(N__14386),
            .I(N__14383));
    Span4Mux_s3_h I__2839 (
            .O(N__14383),
            .I(N__14380));
    Odrv4 I__2838 (
            .O(N__14380),
            .I(\Lab_UT.scctrl.g0_14_mb_rn_0 ));
    CascadeMux I__2837 (
            .O(N__14377),
            .I(\Lab_UT.scctrl.g0_0_i_1_cascade_ ));
    InMux I__2836 (
            .O(N__14374),
            .I(N__14371));
    LocalMux I__2835 (
            .O(N__14371),
            .I(\Lab_UT.scctrl.N_7_2 ));
    InMux I__2834 (
            .O(N__14368),
            .I(N__14365));
    LocalMux I__2833 (
            .O(N__14365),
            .I(N__14362));
    Odrv4 I__2832 (
            .O(N__14362),
            .I(\Lab_UT.scctrl.state_i_3_fast_2 ));
    InMux I__2831 (
            .O(N__14359),
            .I(N__14356));
    LocalMux I__2830 (
            .O(N__14356),
            .I(N__14353));
    Span4Mux_h I__2829 (
            .O(N__14353),
            .I(N__14350));
    Odrv4 I__2828 (
            .O(N__14350),
            .I(\Lab_UT.scctrl.next_state_1_0_a5_0_0_3 ));
    InMux I__2827 (
            .O(N__14347),
            .I(N__14343));
    InMux I__2826 (
            .O(N__14346),
            .I(N__14340));
    LocalMux I__2825 (
            .O(N__14343),
            .I(\Lab_UT.scctrl.g0_i_4 ));
    LocalMux I__2824 (
            .O(N__14340),
            .I(\Lab_UT.scctrl.g0_i_4 ));
    InMux I__2823 (
            .O(N__14335),
            .I(N__14332));
    LocalMux I__2822 (
            .O(N__14332),
            .I(N__14328));
    InMux I__2821 (
            .O(N__14331),
            .I(N__14325));
    Odrv4 I__2820 (
            .O(N__14328),
            .I(\Lab_UT.scctrl.N_10 ));
    LocalMux I__2819 (
            .O(N__14325),
            .I(\Lab_UT.scctrl.N_10 ));
    CascadeMux I__2818 (
            .O(N__14320),
            .I(\Lab_UT.scctrl.G_23_0_a9_4_2_cascade_ ));
    InMux I__2817 (
            .O(N__14317),
            .I(N__14314));
    LocalMux I__2816 (
            .O(N__14314),
            .I(\Lab_UT.scctrl.G_23_0_3 ));
    InMux I__2815 (
            .O(N__14311),
            .I(N__14305));
    InMux I__2814 (
            .O(N__14310),
            .I(N__14305));
    LocalMux I__2813 (
            .O(N__14305),
            .I(\Lab_UT.scctrl.G_23_0_a9_3_1 ));
    InMux I__2812 (
            .O(N__14302),
            .I(N__14296));
    InMux I__2811 (
            .O(N__14301),
            .I(N__14296));
    LocalMux I__2810 (
            .O(N__14296),
            .I(\Lab_UT.scctrl.G_23_0_4 ));
    CascadeMux I__2809 (
            .O(N__14293),
            .I(\Lab_UT.scctrl.G_23_0_3_cascade_ ));
    InMux I__2808 (
            .O(N__14290),
            .I(N__14286));
    InMux I__2807 (
            .O(N__14289),
            .I(N__14283));
    LocalMux I__2806 (
            .O(N__14286),
            .I(\Lab_UT.scctrl.N_3ctr ));
    LocalMux I__2805 (
            .O(N__14283),
            .I(\Lab_UT.scctrl.N_3ctr ));
    CascadeMux I__2804 (
            .O(N__14278),
            .I(N__14275));
    InMux I__2803 (
            .O(N__14275),
            .I(N__14272));
    LocalMux I__2802 (
            .O(N__14272),
            .I(\Lab_UT.scctrl.g0_i_a7_2_0 ));
    CascadeMux I__2801 (
            .O(N__14269),
            .I(N__14266));
    InMux I__2800 (
            .O(N__14266),
            .I(N__14263));
    LocalMux I__2799 (
            .O(N__14263),
            .I(N__14260));
    Span4Mux_v I__2798 (
            .O(N__14260),
            .I(N__14257));
    Odrv4 I__2797 (
            .O(N__14257),
            .I(\Lab_UT.scctrl.next_state_1_i_a5_4_0_0 ));
    InMux I__2796 (
            .O(N__14254),
            .I(N__14251));
    LocalMux I__2795 (
            .O(N__14251),
            .I(\Lab_UT.scctrl.N_8_0 ));
    InMux I__2794 (
            .O(N__14248),
            .I(N__14245));
    LocalMux I__2793 (
            .O(N__14245),
            .I(\Lab_UT.scctrl.g0_i_a9_1 ));
    CascadeMux I__2792 (
            .O(N__14242),
            .I(\Lab_UT.scctrl.N_12_cascade_ ));
    InMux I__2791 (
            .O(N__14239),
            .I(N__14236));
    LocalMux I__2790 (
            .O(N__14236),
            .I(\Lab_UT.scctrl.g0_i_2 ));
    CascadeMux I__2789 (
            .O(N__14233),
            .I(N__14230));
    InMux I__2788 (
            .O(N__14230),
            .I(N__14227));
    LocalMux I__2787 (
            .O(N__14227),
            .I(N__14224));
    Odrv4 I__2786 (
            .O(N__14224),
            .I(\Lab_UT.scctrl.G_23_0_a9_0_0 ));
    CascadeMux I__2785 (
            .O(N__14221),
            .I(\Lab_UT.scctrl.g0_i_a10_2_1_cascade_ ));
    InMux I__2784 (
            .O(N__14218),
            .I(N__14215));
    LocalMux I__2783 (
            .O(N__14215),
            .I(\Lab_UT.scctrl.G_23_0_2 ));
    InMux I__2782 (
            .O(N__14212),
            .I(N__14209));
    LocalMux I__2781 (
            .O(N__14209),
            .I(\Lab_UT.scctrl.N_2ctr ));
    InMux I__2780 (
            .O(N__14206),
            .I(N__14203));
    LocalMux I__2779 (
            .O(N__14203),
            .I(\Lab_UT.scctrl.g0_i_0 ));
    InMux I__2778 (
            .O(N__14200),
            .I(N__14195));
    InMux I__2777 (
            .O(N__14199),
            .I(N__14189));
    InMux I__2776 (
            .O(N__14198),
            .I(N__14189));
    LocalMux I__2775 (
            .O(N__14195),
            .I(N__14186));
    InMux I__2774 (
            .O(N__14194),
            .I(N__14183));
    LocalMux I__2773 (
            .O(N__14189),
            .I(\Lab_UT.state_ret_13_RNIHUNI41_0 ));
    Odrv4 I__2772 (
            .O(N__14186),
            .I(\Lab_UT.state_ret_13_RNIHUNI41_0 ));
    LocalMux I__2771 (
            .O(N__14183),
            .I(\Lab_UT.state_ret_13_RNIHUNI41_0 ));
    CascadeMux I__2770 (
            .O(N__14176),
            .I(\Lab_UT.state_ret_13_RNIHUNI41_0_cascade_ ));
    InMux I__2769 (
            .O(N__14173),
            .I(N__14170));
    LocalMux I__2768 (
            .O(N__14170),
            .I(N__14166));
    InMux I__2767 (
            .O(N__14169),
            .I(N__14163));
    Span4Mux_h I__2766 (
            .O(N__14166),
            .I(N__14160));
    LocalMux I__2765 (
            .O(N__14163),
            .I(\Lab_UT.scdp.key1_2 ));
    Odrv4 I__2764 (
            .O(N__14160),
            .I(\Lab_UT.scdp.key1_2 ));
    CascadeMux I__2763 (
            .O(N__14155),
            .I(N__14150));
    InMux I__2762 (
            .O(N__14154),
            .I(N__14147));
    InMux I__2761 (
            .O(N__14153),
            .I(N__14141));
    InMux I__2760 (
            .O(N__14150),
            .I(N__14141));
    LocalMux I__2759 (
            .O(N__14147),
            .I(N__14138));
    InMux I__2758 (
            .O(N__14146),
            .I(N__14135));
    LocalMux I__2757 (
            .O(N__14141),
            .I(N__14132));
    Span12Mux_s5_v I__2756 (
            .O(N__14138),
            .I(N__14129));
    LocalMux I__2755 (
            .O(N__14135),
            .I(N__14124));
    Span12Mux_s10_v I__2754 (
            .O(N__14132),
            .I(N__14124));
    Odrv12 I__2753 (
            .O(N__14129),
            .I(\Lab_UT.sccDecrypt_0 ));
    Odrv12 I__2752 (
            .O(N__14124),
            .I(\Lab_UT.sccDecrypt_0 ));
    InMux I__2751 (
            .O(N__14119),
            .I(N__14114));
    InMux I__2750 (
            .O(N__14118),
            .I(N__14109));
    InMux I__2749 (
            .O(N__14117),
            .I(N__14109));
    LocalMux I__2748 (
            .O(N__14114),
            .I(\Lab_UT.state_ret_12_RNIMJCP8_0 ));
    LocalMux I__2747 (
            .O(N__14109),
            .I(\Lab_UT.state_ret_12_RNIMJCP8_0 ));
    CascadeMux I__2746 (
            .O(N__14104),
            .I(\Lab_UT.sccDnibble2En_cascade_ ));
    InMux I__2745 (
            .O(N__14101),
            .I(N__14098));
    LocalMux I__2744 (
            .O(N__14098),
            .I(N__14095));
    Span4Mux_h I__2743 (
            .O(N__14095),
            .I(N__14091));
    InMux I__2742 (
            .O(N__14094),
            .I(N__14088));
    Span4Mux_v I__2741 (
            .O(N__14091),
            .I(N__14083));
    LocalMux I__2740 (
            .O(N__14088),
            .I(N__14080));
    InMux I__2739 (
            .O(N__14087),
            .I(N__14077));
    IoInMux I__2738 (
            .O(N__14086),
            .I(N__14074));
    Span4Mux_v I__2737 (
            .O(N__14083),
            .I(N__14069));
    Span4Mux_h I__2736 (
            .O(N__14080),
            .I(N__14069));
    LocalMux I__2735 (
            .O(N__14077),
            .I(N__14066));
    LocalMux I__2734 (
            .O(N__14074),
            .I(N__14063));
    Span4Mux_h I__2733 (
            .O(N__14069),
            .I(N__14060));
    Span4Mux_h I__2732 (
            .O(N__14066),
            .I(N__14057));
    Span4Mux_s1_h I__2731 (
            .O(N__14063),
            .I(N__14054));
    Odrv4 I__2730 (
            .O(N__14060),
            .I(resetGen_rst_0_iso));
    Odrv4 I__2729 (
            .O(N__14057),
            .I(resetGen_rst_0_iso));
    Odrv4 I__2728 (
            .O(N__14054),
            .I(resetGen_rst_0_iso));
    CEMux I__2727 (
            .O(N__14047),
            .I(N__14044));
    LocalMux I__2726 (
            .O(N__14044),
            .I(\Lab_UT.scdp.u1.sccDnibble2En_0 ));
    InMux I__2725 (
            .O(N__14041),
            .I(N__14037));
    InMux I__2724 (
            .O(N__14040),
            .I(N__14034));
    LocalMux I__2723 (
            .O(N__14037),
            .I(N__14031));
    LocalMux I__2722 (
            .O(N__14034),
            .I(N__14028));
    Span4Mux_s2_v I__2721 (
            .O(N__14031),
            .I(N__14023));
    Span4Mux_h I__2720 (
            .O(N__14028),
            .I(N__14023));
    Odrv4 I__2719 (
            .O(N__14023),
            .I(\Lab_UT.scdp.N_37 ));
    InMux I__2718 (
            .O(N__14020),
            .I(N__14014));
    InMux I__2717 (
            .O(N__14019),
            .I(N__14014));
    LocalMux I__2716 (
            .O(N__14014),
            .I(N__14010));
    InMux I__2715 (
            .O(N__14013),
            .I(N__14007));
    Odrv4 I__2714 (
            .O(N__14010),
            .I(\Lab_UT.sccDnibble2En ));
    LocalMux I__2713 (
            .O(N__14007),
            .I(\Lab_UT.sccDnibble2En ));
    InMux I__2712 (
            .O(N__14002),
            .I(N__13998));
    CascadeMux I__2711 (
            .O(N__14001),
            .I(N__13995));
    LocalMux I__2710 (
            .O(N__13998),
            .I(N__13992));
    InMux I__2709 (
            .O(N__13995),
            .I(N__13989));
    Span4Mux_h I__2708 (
            .O(N__13992),
            .I(N__13985));
    LocalMux I__2707 (
            .O(N__13989),
            .I(N__13982));
    InMux I__2706 (
            .O(N__13988),
            .I(N__13979));
    Span4Mux_v I__2705 (
            .O(N__13985),
            .I(N__13976));
    Span4Mux_h I__2704 (
            .O(N__13982),
            .I(N__13973));
    LocalMux I__2703 (
            .O(N__13979),
            .I(\Lab_UT.scdp.byteToDecrypt_1 ));
    Odrv4 I__2702 (
            .O(N__13976),
            .I(\Lab_UT.scdp.byteToDecrypt_1 ));
    Odrv4 I__2701 (
            .O(N__13973),
            .I(\Lab_UT.scdp.byteToDecrypt_1 ));
    IoInMux I__2700 (
            .O(N__13966),
            .I(N__13960));
    CascadeMux I__2699 (
            .O(N__13965),
            .I(N__13957));
    InMux I__2698 (
            .O(N__13964),
            .I(N__13954));
    InMux I__2697 (
            .O(N__13963),
            .I(N__13951));
    LocalMux I__2696 (
            .O(N__13960),
            .I(N__13948));
    InMux I__2695 (
            .O(N__13957),
            .I(N__13945));
    LocalMux I__2694 (
            .O(N__13954),
            .I(N__13942));
    LocalMux I__2693 (
            .O(N__13951),
            .I(N__13939));
    IoSpan4Mux I__2692 (
            .O(N__13948),
            .I(N__13936));
    LocalMux I__2691 (
            .O(N__13945),
            .I(N__13933));
    Span4Mux_v I__2690 (
            .O(N__13942),
            .I(N__13930));
    Span4Mux_h I__2689 (
            .O(N__13939),
            .I(N__13923));
    Span4Mux_s1_v I__2688 (
            .O(N__13936),
            .I(N__13923));
    Span4Mux_v I__2687 (
            .O(N__13933),
            .I(N__13923));
    Odrv4 I__2686 (
            .O(N__13930),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2685 (
            .O(N__13923),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__2684 (
            .O(N__13918),
            .I(\Lab_UT.scctrl.g0_i_a9_0_1_cascade_ ));
    InMux I__2683 (
            .O(N__13915),
            .I(N__13912));
    LocalMux I__2682 (
            .O(N__13912),
            .I(N__13908));
    InMux I__2681 (
            .O(N__13911),
            .I(N__13905));
    Odrv4 I__2680 (
            .O(N__13908),
            .I(\Lab_UT.scctrl.next_state77_2 ));
    LocalMux I__2679 (
            .O(N__13905),
            .I(\Lab_UT.scctrl.next_state77_2 ));
    InMux I__2678 (
            .O(N__13900),
            .I(N__13897));
    LocalMux I__2677 (
            .O(N__13897),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz_4 ));
    InMux I__2676 (
            .O(N__13894),
            .I(N__13891));
    LocalMux I__2675 (
            .O(N__13891),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz ));
    CascadeMux I__2674 (
            .O(N__13888),
            .I(N__13885));
    InMux I__2673 (
            .O(N__13885),
            .I(N__13879));
    InMux I__2672 (
            .O(N__13884),
            .I(N__13879));
    LocalMux I__2671 (
            .O(N__13879),
            .I(N__13876));
    Odrv12 I__2670 (
            .O(N__13876),
            .I(\Lab_UT.scctrl.next_state76 ));
    InMux I__2669 (
            .O(N__13873),
            .I(N__13870));
    LocalMux I__2668 (
            .O(N__13870),
            .I(N__13866));
    InMux I__2667 (
            .O(N__13869),
            .I(N__13863));
    Span4Mux_h I__2666 (
            .O(N__13866),
            .I(N__13860));
    LocalMux I__2665 (
            .O(N__13863),
            .I(\Lab_UT.scdp.key2_3 ));
    Odrv4 I__2664 (
            .O(N__13860),
            .I(\Lab_UT.scdp.key2_3 ));
    InMux I__2663 (
            .O(N__13855),
            .I(N__13852));
    LocalMux I__2662 (
            .O(N__13852),
            .I(N__13848));
    InMux I__2661 (
            .O(N__13851),
            .I(N__13845));
    Span4Mux_h I__2660 (
            .O(N__13848),
            .I(N__13842));
    LocalMux I__2659 (
            .O(N__13845),
            .I(\Lab_UT.scdp.key2_6 ));
    Odrv4 I__2658 (
            .O(N__13842),
            .I(\Lab_UT.scdp.key2_6 ));
    InMux I__2657 (
            .O(N__13837),
            .I(N__13831));
    InMux I__2656 (
            .O(N__13836),
            .I(N__13828));
    InMux I__2655 (
            .O(N__13835),
            .I(N__13823));
    InMux I__2654 (
            .O(N__13834),
            .I(N__13823));
    LocalMux I__2653 (
            .O(N__13831),
            .I(\Lab_UT.state_ret_14_RNI416G41_0 ));
    LocalMux I__2652 (
            .O(N__13828),
            .I(\Lab_UT.state_ret_14_RNI416G41_0 ));
    LocalMux I__2651 (
            .O(N__13823),
            .I(\Lab_UT.state_ret_14_RNI416G41_0 ));
    InMux I__2650 (
            .O(N__13816),
            .I(N__13812));
    CascadeMux I__2649 (
            .O(N__13815),
            .I(N__13809));
    LocalMux I__2648 (
            .O(N__13812),
            .I(N__13806));
    InMux I__2647 (
            .O(N__13809),
            .I(N__13803));
    Span4Mux_h I__2646 (
            .O(N__13806),
            .I(N__13800));
    LocalMux I__2645 (
            .O(N__13803),
            .I(\Lab_UT.scdp.key3_6 ));
    Odrv4 I__2644 (
            .O(N__13800),
            .I(\Lab_UT.scdp.key3_6 ));
    CascadeMux I__2643 (
            .O(N__13795),
            .I(N__13792));
    InMux I__2642 (
            .O(N__13792),
            .I(N__13788));
    CascadeMux I__2641 (
            .O(N__13791),
            .I(N__13785));
    LocalMux I__2640 (
            .O(N__13788),
            .I(N__13782));
    InMux I__2639 (
            .O(N__13785),
            .I(N__13779));
    Span4Mux_v I__2638 (
            .O(N__13782),
            .I(N__13776));
    LocalMux I__2637 (
            .O(N__13779),
            .I(\Lab_UT.scdp.key3_2 ));
    Odrv4 I__2636 (
            .O(N__13776),
            .I(\Lab_UT.scdp.key3_2 ));
    InMux I__2635 (
            .O(N__13771),
            .I(N__13764));
    InMux I__2634 (
            .O(N__13770),
            .I(N__13759));
    InMux I__2633 (
            .O(N__13769),
            .I(N__13759));
    InMux I__2632 (
            .O(N__13768),
            .I(N__13754));
    InMux I__2631 (
            .O(N__13767),
            .I(N__13754));
    LocalMux I__2630 (
            .O(N__13764),
            .I(\Lab_UT.state_2_RNI44QH41_0_2 ));
    LocalMux I__2629 (
            .O(N__13759),
            .I(\Lab_UT.state_2_RNI44QH41_0_2 ));
    LocalMux I__2628 (
            .O(N__13754),
            .I(\Lab_UT.state_2_RNI44QH41_0_2 ));
    InMux I__2627 (
            .O(N__13747),
            .I(N__13744));
    LocalMux I__2626 (
            .O(N__13744),
            .I(N__13741));
    Span4Mux_v I__2625 (
            .O(N__13741),
            .I(N__13737));
    InMux I__2624 (
            .O(N__13740),
            .I(N__13734));
    Span4Mux_s2_v I__2623 (
            .O(N__13737),
            .I(N__13731));
    LocalMux I__2622 (
            .O(N__13734),
            .I(\Lab_UT.scdp.key2_7 ));
    Odrv4 I__2621 (
            .O(N__13731),
            .I(\Lab_UT.scdp.key2_7 ));
    InMux I__2620 (
            .O(N__13726),
            .I(N__13719));
    InMux I__2619 (
            .O(N__13725),
            .I(N__13714));
    InMux I__2618 (
            .O(N__13724),
            .I(N__13714));
    InMux I__2617 (
            .O(N__13723),
            .I(N__13711));
    InMux I__2616 (
            .O(N__13722),
            .I(N__13708));
    LocalMux I__2615 (
            .O(N__13719),
            .I(\Lab_UT.state_2_RNIF0RJ41_0_2 ));
    LocalMux I__2614 (
            .O(N__13714),
            .I(\Lab_UT.state_2_RNIF0RJ41_0_2 ));
    LocalMux I__2613 (
            .O(N__13711),
            .I(\Lab_UT.state_2_RNIF0RJ41_0_2 ));
    LocalMux I__2612 (
            .O(N__13708),
            .I(\Lab_UT.state_2_RNIF0RJ41_0_2 ));
    InMux I__2611 (
            .O(N__13699),
            .I(N__13696));
    LocalMux I__2610 (
            .O(N__13696),
            .I(N__13692));
    InMux I__2609 (
            .O(N__13695),
            .I(N__13689));
    Span4Mux_h I__2608 (
            .O(N__13692),
            .I(N__13686));
    LocalMux I__2607 (
            .O(N__13689),
            .I(\Lab_UT.scdp.key3_3 ));
    Odrv4 I__2606 (
            .O(N__13686),
            .I(\Lab_UT.scdp.key3_3 ));
    InMux I__2605 (
            .O(N__13681),
            .I(N__13677));
    InMux I__2604 (
            .O(N__13680),
            .I(N__13674));
    LocalMux I__2603 (
            .O(N__13677),
            .I(\Lab_UT.scdp.key0_0 ));
    LocalMux I__2602 (
            .O(N__13674),
            .I(\Lab_UT.scdp.key0_0 ));
    CascadeMux I__2601 (
            .O(N__13669),
            .I(N__13666));
    InMux I__2600 (
            .O(N__13666),
            .I(N__13662));
    InMux I__2599 (
            .O(N__13665),
            .I(N__13659));
    LocalMux I__2598 (
            .O(N__13662),
            .I(\Lab_UT.scdp.key0_2 ));
    LocalMux I__2597 (
            .O(N__13659),
            .I(\Lab_UT.scdp.key0_2 ));
    InMux I__2596 (
            .O(N__13654),
            .I(N__13650));
    InMux I__2595 (
            .O(N__13653),
            .I(N__13647));
    LocalMux I__2594 (
            .O(N__13650),
            .I(N__13644));
    LocalMux I__2593 (
            .O(N__13647),
            .I(\Lab_UT.scdp.key1_4 ));
    Odrv4 I__2592 (
            .O(N__13644),
            .I(\Lab_UT.scdp.key1_4 ));
    InMux I__2591 (
            .O(N__13639),
            .I(N__13632));
    InMux I__2590 (
            .O(N__13638),
            .I(N__13629));
    InMux I__2589 (
            .O(N__13637),
            .I(N__13626));
    InMux I__2588 (
            .O(N__13636),
            .I(N__13621));
    InMux I__2587 (
            .O(N__13635),
            .I(N__13621));
    LocalMux I__2586 (
            .O(N__13632),
            .I(N__13618));
    LocalMux I__2585 (
            .O(N__13629),
            .I(\Lab_UT.state_ret_13_RNIQ72741_0 ));
    LocalMux I__2584 (
            .O(N__13626),
            .I(\Lab_UT.state_ret_13_RNIQ72741_0 ));
    LocalMux I__2583 (
            .O(N__13621),
            .I(\Lab_UT.state_ret_13_RNIQ72741_0 ));
    Odrv4 I__2582 (
            .O(N__13618),
            .I(\Lab_UT.state_ret_13_RNIQ72741_0 ));
    InMux I__2581 (
            .O(N__13609),
            .I(N__13606));
    LocalMux I__2580 (
            .O(N__13606),
            .I(N__13603));
    Span4Mux_h I__2579 (
            .O(N__13603),
            .I(N__13599));
    InMux I__2578 (
            .O(N__13602),
            .I(N__13596));
    Span4Mux_h I__2577 (
            .O(N__13599),
            .I(N__13593));
    LocalMux I__2576 (
            .O(N__13596),
            .I(\Lab_UT.scdp.key1_6 ));
    Odrv4 I__2575 (
            .O(N__13593),
            .I(\Lab_UT.scdp.key1_6 ));
    CascadeMux I__2574 (
            .O(N__13588),
            .I(\Lab_UT.scctrl.next_state77_cascade_ ));
    InMux I__2573 (
            .O(N__13585),
            .I(N__13580));
    InMux I__2572 (
            .O(N__13584),
            .I(N__13575));
    InMux I__2571 (
            .O(N__13583),
            .I(N__13575));
    LocalMux I__2570 (
            .O(N__13580),
            .I(N__13572));
    LocalMux I__2569 (
            .O(N__13575),
            .I(\Lab_UT.scctrl.next_state_3_sqmuxa ));
    Odrv4 I__2568 (
            .O(N__13572),
            .I(\Lab_UT.scctrl.next_state_3_sqmuxa ));
    CascadeMux I__2567 (
            .O(N__13567),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_0_cascade_ ));
    InMux I__2566 (
            .O(N__13564),
            .I(N__13561));
    LocalMux I__2565 (
            .O(N__13561),
            .I(\Lab_UT.scctrl.next_state77 ));
    CascadeMux I__2564 (
            .O(N__13558),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_cascade_ ));
    CascadeMux I__2563 (
            .O(N__13555),
            .I(\Lab_UT.scctrl.g0_i_a9_3_4_cascade_ ));
    InMux I__2562 (
            .O(N__13552),
            .I(N__13549));
    LocalMux I__2561 (
            .O(N__13549),
            .I(N__13546));
    Span4Mux_s3_v I__2560 (
            .O(N__13546),
            .I(N__13543));
    Span4Mux_v I__2559 (
            .O(N__13543),
            .I(N__13540));
    Odrv4 I__2558 (
            .O(N__13540),
            .I(\Lab_UT.scctrl.g0_i_a9_3_5 ));
    CascadeMux I__2557 (
            .O(N__13537),
            .I(\Lab_UT.scctrl.next_state_1_0_a5_2_out_cascade_ ));
    InMux I__2556 (
            .O(N__13534),
            .I(N__13531));
    LocalMux I__2555 (
            .O(N__13531),
            .I(\Lab_UT.scctrl.N_222_1 ));
    InMux I__2554 (
            .O(N__13528),
            .I(N__13525));
    LocalMux I__2553 (
            .O(N__13525),
            .I(N__13522));
    Odrv4 I__2552 (
            .O(N__13522),
            .I(\Lab_UT.scctrl.next_state_3_sqmuxa_0 ));
    InMux I__2551 (
            .O(N__13519),
            .I(N__13516));
    LocalMux I__2550 (
            .O(N__13516),
            .I(N__13513));
    Odrv12 I__2549 (
            .O(N__13513),
            .I(\Lab_UT.scdp.a2b.g1_1_a3_0Z0Z_0 ));
    CascadeMux I__2548 (
            .O(N__13510),
            .I(N__13506));
    InMux I__2547 (
            .O(N__13509),
            .I(N__13503));
    InMux I__2546 (
            .O(N__13506),
            .I(N__13500));
    LocalMux I__2545 (
            .O(N__13503),
            .I(buart__rx_shifter_ret_1_fast));
    LocalMux I__2544 (
            .O(N__13500),
            .I(buart__rx_shifter_ret_1_fast));
    CascadeMux I__2543 (
            .O(N__13495),
            .I(N__13492));
    InMux I__2542 (
            .O(N__13492),
            .I(N__13489));
    LocalMux I__2541 (
            .O(N__13489),
            .I(N__13486));
    Odrv12 I__2540 (
            .O(N__13486),
            .I(\Lab_UT.scctrl.g0_i_o9_0Z0Z_2 ));
    InMux I__2539 (
            .O(N__13483),
            .I(N__13477));
    InMux I__2538 (
            .O(N__13482),
            .I(N__13477));
    LocalMux I__2537 (
            .O(N__13477),
            .I(\Lab_UT.dk.un4_de_hexZ0Z_1 ));
    InMux I__2536 (
            .O(N__13474),
            .I(N__13470));
    CascadeMux I__2535 (
            .O(N__13473),
            .I(N__13465));
    LocalMux I__2534 (
            .O(N__13470),
            .I(N__13461));
    InMux I__2533 (
            .O(N__13469),
            .I(N__13456));
    InMux I__2532 (
            .O(N__13468),
            .I(N__13456));
    InMux I__2531 (
            .O(N__13465),
            .I(N__13453));
    InMux I__2530 (
            .O(N__13464),
            .I(N__13450));
    Span4Mux_h I__2529 (
            .O(N__13461),
            .I(N__13447));
    LocalMux I__2528 (
            .O(N__13456),
            .I(bu_rx_data_i_3_4));
    LocalMux I__2527 (
            .O(N__13453),
            .I(bu_rx_data_i_3_4));
    LocalMux I__2526 (
            .O(N__13450),
            .I(bu_rx_data_i_3_4));
    Odrv4 I__2525 (
            .O(N__13447),
            .I(bu_rx_data_i_3_4));
    InMux I__2524 (
            .O(N__13438),
            .I(N__13434));
    InMux I__2523 (
            .O(N__13437),
            .I(N__13430));
    LocalMux I__2522 (
            .O(N__13434),
            .I(N__13427));
    InMux I__2521 (
            .O(N__13433),
            .I(N__13424));
    LocalMux I__2520 (
            .O(N__13430),
            .I(N__13421));
    Span4Mux_s3_h I__2519 (
            .O(N__13427),
            .I(N__13418));
    LocalMux I__2518 (
            .O(N__13424),
            .I(N__13413));
    Span4Mux_s3_h I__2517 (
            .O(N__13421),
            .I(N__13413));
    Span4Mux_h I__2516 (
            .O(N__13418),
            .I(N__13401));
    Span4Mux_h I__2515 (
            .O(N__13413),
            .I(N__13401));
    InMux I__2514 (
            .O(N__13412),
            .I(N__13396));
    InMux I__2513 (
            .O(N__13411),
            .I(N__13396));
    InMux I__2512 (
            .O(N__13410),
            .I(N__13385));
    InMux I__2511 (
            .O(N__13409),
            .I(N__13385));
    InMux I__2510 (
            .O(N__13408),
            .I(N__13385));
    InMux I__2509 (
            .O(N__13407),
            .I(N__13385));
    InMux I__2508 (
            .O(N__13406),
            .I(N__13385));
    Odrv4 I__2507 (
            .O(N__13401),
            .I(bu_rx_data_5));
    LocalMux I__2506 (
            .O(N__13396),
            .I(bu_rx_data_5));
    LocalMux I__2505 (
            .O(N__13385),
            .I(bu_rx_data_5));
    InMux I__2504 (
            .O(N__13378),
            .I(N__13370));
    InMux I__2503 (
            .O(N__13377),
            .I(N__13365));
    InMux I__2502 (
            .O(N__13376),
            .I(N__13365));
    InMux I__2501 (
            .O(N__13375),
            .I(N__13358));
    InMux I__2500 (
            .O(N__13374),
            .I(N__13358));
    InMux I__2499 (
            .O(N__13373),
            .I(N__13358));
    LocalMux I__2498 (
            .O(N__13370),
            .I(N__13354));
    LocalMux I__2497 (
            .O(N__13365),
            .I(N__13351));
    LocalMux I__2496 (
            .O(N__13358),
            .I(N__13346));
    InMux I__2495 (
            .O(N__13357),
            .I(N__13343));
    Span12Mux_s6_v I__2494 (
            .O(N__13354),
            .I(N__13338));
    Span12Mux_s9_v I__2493 (
            .O(N__13351),
            .I(N__13338));
    InMux I__2492 (
            .O(N__13350),
            .I(N__13333));
    InMux I__2491 (
            .O(N__13349),
            .I(N__13333));
    Odrv4 I__2490 (
            .O(N__13346),
            .I(bu_rx_data_4));
    LocalMux I__2489 (
            .O(N__13343),
            .I(bu_rx_data_4));
    Odrv12 I__2488 (
            .O(N__13338),
            .I(bu_rx_data_4));
    LocalMux I__2487 (
            .O(N__13333),
            .I(bu_rx_data_4));
    CascadeMux I__2486 (
            .O(N__13324),
            .I(N__13319));
    CascadeMux I__2485 (
            .O(N__13323),
            .I(N__13315));
    CascadeMux I__2484 (
            .O(N__13322),
            .I(N__13312));
    InMux I__2483 (
            .O(N__13319),
            .I(N__13309));
    InMux I__2482 (
            .O(N__13318),
            .I(N__13306));
    InMux I__2481 (
            .O(N__13315),
            .I(N__13300));
    InMux I__2480 (
            .O(N__13312),
            .I(N__13300));
    LocalMux I__2479 (
            .O(N__13309),
            .I(N__13297));
    LocalMux I__2478 (
            .O(N__13306),
            .I(N__13294));
    InMux I__2477 (
            .O(N__13305),
            .I(N__13291));
    LocalMux I__2476 (
            .O(N__13300),
            .I(N__13288));
    Odrv4 I__2475 (
            .O(N__13297),
            .I(bu_rx_data_i_2_6));
    Odrv12 I__2474 (
            .O(N__13294),
            .I(bu_rx_data_i_2_6));
    LocalMux I__2473 (
            .O(N__13291),
            .I(bu_rx_data_i_2_6));
    Odrv4 I__2472 (
            .O(N__13288),
            .I(bu_rx_data_i_2_6));
    InMux I__2471 (
            .O(N__13279),
            .I(N__13275));
    InMux I__2470 (
            .O(N__13278),
            .I(N__13272));
    LocalMux I__2469 (
            .O(N__13275),
            .I(\Lab_UT.un1_de_hex_2 ));
    LocalMux I__2468 (
            .O(N__13272),
            .I(\Lab_UT.un1_de_hex_2 ));
    CascadeMux I__2467 (
            .O(N__13267),
            .I(\Lab_UT.un1_de_hex_2_cascade_ ));
    InMux I__2466 (
            .O(N__13264),
            .I(N__13261));
    LocalMux I__2465 (
            .O(N__13261),
            .I(\Lab_UT.scctrl.N_9_0 ));
    InMux I__2464 (
            .O(N__13258),
            .I(N__13255));
    LocalMux I__2463 (
            .O(N__13255),
            .I(bu_rx_data_fast_0));
    InMux I__2462 (
            .O(N__13252),
            .I(N__13247));
    InMux I__2461 (
            .O(N__13251),
            .I(N__13244));
    InMux I__2460 (
            .O(N__13250),
            .I(N__13241));
    LocalMux I__2459 (
            .O(N__13247),
            .I(N__13238));
    LocalMux I__2458 (
            .O(N__13244),
            .I(buart__rx_shifter_0_fast_3));
    LocalMux I__2457 (
            .O(N__13241),
            .I(buart__rx_shifter_0_fast_3));
    Odrv4 I__2456 (
            .O(N__13238),
            .I(buart__rx_shifter_0_fast_3));
    CascadeMux I__2455 (
            .O(N__13231),
            .I(\Lab_UT.dk.un7_de_hex_xZ0Z0_cascade_ ));
    CascadeMux I__2454 (
            .O(N__13228),
            .I(\Lab_UT.dk.un7_de_hex_0_cascade_ ));
    InMux I__2453 (
            .O(N__13225),
            .I(N__13222));
    LocalMux I__2452 (
            .O(N__13222),
            .I(\Lab_UT.dk.un7_de_hex_0 ));
    CascadeMux I__2451 (
            .O(N__13219),
            .I(\Lab_UT.un4_de_hex_cascade_ ));
    InMux I__2450 (
            .O(N__13216),
            .I(N__13213));
    LocalMux I__2449 (
            .O(N__13213),
            .I(buart__rx_shifter_0_fast_1));
    CascadeMux I__2448 (
            .O(N__13210),
            .I(\Lab_UT.scctrl.EmsLoaded_cascade_ ));
    CascadeMux I__2447 (
            .O(N__13207),
            .I(\Lab_UT.sccElsBitsLd_cascade_ ));
    CEMux I__2446 (
            .O(N__13204),
            .I(N__13201));
    LocalMux I__2445 (
            .O(N__13201),
            .I(N__13197));
    CEMux I__2444 (
            .O(N__13200),
            .I(N__13194));
    Span4Mux_v I__2443 (
            .O(N__13197),
            .I(N__13189));
    LocalMux I__2442 (
            .O(N__13194),
            .I(N__13189));
    Span4Mux_v I__2441 (
            .O(N__13189),
            .I(N__13186));
    Odrv4 I__2440 (
            .O(N__13186),
            .I(\Lab_UT.scdp.sccElsBitsLd_0 ));
    InMux I__2439 (
            .O(N__13183),
            .I(N__13174));
    InMux I__2438 (
            .O(N__13182),
            .I(N__13174));
    InMux I__2437 (
            .O(N__13181),
            .I(N__13174));
    LocalMux I__2436 (
            .O(N__13174),
            .I(N__13171));
    Span4Mux_v I__2435 (
            .O(N__13171),
            .I(N__13167));
    InMux I__2434 (
            .O(N__13170),
            .I(N__13164));
    Span4Mux_v I__2433 (
            .O(N__13167),
            .I(N__13161));
    LocalMux I__2432 (
            .O(N__13164),
            .I(\Lab_UT.sccElsBitsLd ));
    Odrv4 I__2431 (
            .O(N__13161),
            .I(\Lab_UT.sccElsBitsLd ));
    CascadeMux I__2430 (
            .O(N__13156),
            .I(N__13153));
    InMux I__2429 (
            .O(N__13153),
            .I(N__13150));
    LocalMux I__2428 (
            .O(N__13150),
            .I(N__13147));
    Span4Mux_v I__2427 (
            .O(N__13147),
            .I(N__13143));
    InMux I__2426 (
            .O(N__13146),
            .I(N__13140));
    Odrv4 I__2425 (
            .O(N__13143),
            .I(\Lab_UT.scdp.lsBitsi.lsBitsD_5 ));
    LocalMux I__2424 (
            .O(N__13140),
            .I(\Lab_UT.scdp.lsBitsi.lsBitsD_5 ));
    CascadeMux I__2423 (
            .O(N__13135),
            .I(Lab_UT_dk_de_cr_12_1_cascade_));
    CascadeMux I__2422 (
            .O(N__13132),
            .I(L4_PrintBuf_cascade_));
    CascadeMux I__2421 (
            .O(N__13129),
            .I(\Lab_UT.sccDnibble1En_cascade_ ));
    CEMux I__2420 (
            .O(N__13126),
            .I(N__13123));
    LocalMux I__2419 (
            .O(N__13123),
            .I(N__13120));
    Span4Mux_v I__2418 (
            .O(N__13120),
            .I(N__13117));
    Odrv4 I__2417 (
            .O(N__13117),
            .I(\Lab_UT.scdp.u0.sccDnibble1En_0 ));
    CascadeMux I__2416 (
            .O(N__13114),
            .I(\Lab_UT.scctrl.next_state_1_sqmuxa_3_0_cascade_ ));
    InMux I__2415 (
            .O(N__13111),
            .I(N__13105));
    InMux I__2414 (
            .O(N__13110),
            .I(N__13105));
    LocalMux I__2413 (
            .O(N__13105),
            .I(N__13102));
    Odrv4 I__2412 (
            .O(N__13102),
            .I(\Lab_UT.scctrl.state_retZ0Z_10 ));
    CascadeMux I__2411 (
            .O(N__13099),
            .I(\Lab_UT.scctrl.next_state_1_sqmuxa_3_cascade_ ));
    CascadeMux I__2410 (
            .O(N__13096),
            .I(N__13092));
    InMux I__2409 (
            .O(N__13095),
            .I(N__13089));
    InMux I__2408 (
            .O(N__13092),
            .I(N__13086));
    LocalMux I__2407 (
            .O(N__13089),
            .I(\Lab_UT.scctrl.nibbleInZ0Z1 ));
    LocalMux I__2406 (
            .O(N__13086),
            .I(\Lab_UT.scctrl.nibbleInZ0Z1 ));
    CEMux I__2405 (
            .O(N__13081),
            .I(N__13078));
    LocalMux I__2404 (
            .O(N__13078),
            .I(N__13075));
    Span4Mux_v I__2403 (
            .O(N__13075),
            .I(N__13072));
    Span4Mux_s2_v I__2402 (
            .O(N__13072),
            .I(N__13069));
    Odrv4 I__2401 (
            .O(N__13069),
            .I(\Lab_UT.scctrl.N_1_0_i ));
    SRMux I__2400 (
            .O(N__13066),
            .I(N__13063));
    LocalMux I__2399 (
            .O(N__13063),
            .I(N__13060));
    Sp12to4 I__2398 (
            .O(N__13060),
            .I(N__13056));
    InMux I__2397 (
            .O(N__13059),
            .I(N__13053));
    Odrv12 I__2396 (
            .O(N__13056),
            .I(\Lab_UT.scctrl.next_state_1_sqmuxa_3 ));
    LocalMux I__2395 (
            .O(N__13053),
            .I(\Lab_UT.scctrl.next_state_1_sqmuxa_3 ));
    InMux I__2394 (
            .O(N__13048),
            .I(N__13045));
    LocalMux I__2393 (
            .O(N__13045),
            .I(N__13041));
    InMux I__2392 (
            .O(N__13044),
            .I(N__13038));
    Span12Mux_s3_v I__2391 (
            .O(N__13041),
            .I(N__13035));
    LocalMux I__2390 (
            .O(N__13038),
            .I(\Lab_UT.scctrl.un6_sccDecrypt ));
    Odrv12 I__2389 (
            .O(N__13035),
            .I(\Lab_UT.scctrl.un6_sccDecrypt ));
    InMux I__2388 (
            .O(N__13030),
            .I(N__13027));
    LocalMux I__2387 (
            .O(N__13027),
            .I(N__13024));
    Odrv4 I__2386 (
            .O(N__13024),
            .I(\Lab_UT.de_bigE ));
    InMux I__2385 (
            .O(N__13021),
            .I(N__13018));
    LocalMux I__2384 (
            .O(N__13018),
            .I(N__13013));
    InMux I__2383 (
            .O(N__13017),
            .I(N__13010));
    InMux I__2382 (
            .O(N__13016),
            .I(N__13007));
    Odrv4 I__2381 (
            .O(N__13013),
            .I(\Lab_UT.scctrl.next_state_1_i_a5_1_0 ));
    LocalMux I__2380 (
            .O(N__13010),
            .I(\Lab_UT.scctrl.next_state_1_i_a5_1_0 ));
    LocalMux I__2379 (
            .O(N__13007),
            .I(\Lab_UT.scctrl.next_state_1_i_a5_1_0 ));
    InMux I__2378 (
            .O(N__13000),
            .I(N__12997));
    LocalMux I__2377 (
            .O(N__12997),
            .I(\Lab_UT.scctrl.EmsLoaded ));
    InMux I__2376 (
            .O(N__12994),
            .I(N__12991));
    LocalMux I__2375 (
            .O(N__12991),
            .I(N__12988));
    Odrv12 I__2374 (
            .O(N__12988),
            .I(\Lab_UT.scctrl.g0_7_1_0 ));
    CascadeMux I__2373 (
            .O(N__12985),
            .I(\Lab_UT.scctrl.g2_0_2_cascade_ ));
    CascadeMux I__2372 (
            .O(N__12982),
            .I(\Lab_UT.scctrl.g0_2_cascade_ ));
    CascadeMux I__2371 (
            .O(N__12979),
            .I(\Lab_UT.scctrl.g0_7_cascade_ ));
    InMux I__2370 (
            .O(N__12976),
            .I(N__12973));
    LocalMux I__2369 (
            .O(N__12973),
            .I(\Lab_UT.scctrl.g1_0 ));
    InMux I__2368 (
            .O(N__12970),
            .I(N__12967));
    LocalMux I__2367 (
            .O(N__12967),
            .I(N__12964));
    Odrv4 I__2366 (
            .O(N__12964),
            .I(\Lab_UT.scctrl.g2_2 ));
    InMux I__2365 (
            .O(N__12961),
            .I(N__12958));
    LocalMux I__2364 (
            .O(N__12958),
            .I(N__12955));
    Odrv4 I__2363 (
            .O(N__12955),
            .I(\Lab_UT.scctrl.g1 ));
    InMux I__2362 (
            .O(N__12952),
            .I(N__12946));
    InMux I__2361 (
            .O(N__12951),
            .I(N__12946));
    LocalMux I__2360 (
            .O(N__12946),
            .I(N__12942));
    InMux I__2359 (
            .O(N__12945),
            .I(N__12939));
    Span4Mux_v I__2358 (
            .O(N__12942),
            .I(N__12936));
    LocalMux I__2357 (
            .O(N__12939),
            .I(N__12933));
    Span4Mux_v I__2356 (
            .O(N__12936),
            .I(N__12930));
    Span4Mux_v I__2355 (
            .O(N__12933),
            .I(N__12927));
    Odrv4 I__2354 (
            .O(N__12930),
            .I(\Lab_UT.sccDnibble1En ));
    Odrv4 I__2353 (
            .O(N__12927),
            .I(\Lab_UT.sccDnibble1En ));
    CascadeMux I__2352 (
            .O(N__12922),
            .I(\Lab_UT.scctrl.next_state_rst_1_0_cascade_ ));
    CascadeMux I__2351 (
            .O(N__12919),
            .I(\Lab_UT.scctrl.un1_state_3_1_reti_cascade_ ));
    CascadeMux I__2350 (
            .O(N__12916),
            .I(N__12913));
    InMux I__2349 (
            .O(N__12913),
            .I(N__12910));
    LocalMux I__2348 (
            .O(N__12910),
            .I(\Lab_UT.de_bigE_0 ));
    InMux I__2347 (
            .O(N__12907),
            .I(N__12903));
    CascadeMux I__2346 (
            .O(N__12906),
            .I(N__12900));
    LocalMux I__2345 (
            .O(N__12903),
            .I(N__12897));
    InMux I__2344 (
            .O(N__12900),
            .I(N__12894));
    Span4Mux_h I__2343 (
            .O(N__12897),
            .I(N__12891));
    LocalMux I__2342 (
            .O(N__12894),
            .I(\Lab_UT.scdp.key3_1 ));
    Odrv4 I__2341 (
            .O(N__12891),
            .I(\Lab_UT.scdp.key3_1 ));
    CascadeMux I__2340 (
            .O(N__12886),
            .I(N__12882));
    CascadeMux I__2339 (
            .O(N__12885),
            .I(N__12879));
    InMux I__2338 (
            .O(N__12882),
            .I(N__12876));
    InMux I__2337 (
            .O(N__12879),
            .I(N__12873));
    LocalMux I__2336 (
            .O(N__12876),
            .I(N__12870));
    LocalMux I__2335 (
            .O(N__12873),
            .I(\Lab_UT.scdp.key1_0 ));
    Odrv4 I__2334 (
            .O(N__12870),
            .I(\Lab_UT.scdp.key1_0 ));
    CascadeMux I__2333 (
            .O(N__12865),
            .I(N__12861));
    CascadeMux I__2332 (
            .O(N__12864),
            .I(N__12858));
    InMux I__2331 (
            .O(N__12861),
            .I(N__12855));
    InMux I__2330 (
            .O(N__12858),
            .I(N__12852));
    LocalMux I__2329 (
            .O(N__12855),
            .I(N__12849));
    LocalMux I__2328 (
            .O(N__12852),
            .I(N__12846));
    Odrv4 I__2327 (
            .O(N__12849),
            .I(\Lab_UT.scdp.key2_4 ));
    Odrv4 I__2326 (
            .O(N__12846),
            .I(\Lab_UT.scdp.key2_4 ));
    InMux I__2325 (
            .O(N__12841),
            .I(N__12838));
    LocalMux I__2324 (
            .O(N__12838),
            .I(N__12834));
    InMux I__2323 (
            .O(N__12837),
            .I(N__12831));
    Span4Mux_h I__2322 (
            .O(N__12834),
            .I(N__12828));
    LocalMux I__2321 (
            .O(N__12831),
            .I(\Lab_UT.scdp.key3_4 ));
    Odrv4 I__2320 (
            .O(N__12828),
            .I(\Lab_UT.scdp.key3_4 ));
    InMux I__2319 (
            .O(N__12823),
            .I(N__12820));
    LocalMux I__2318 (
            .O(N__12820),
            .I(N__12816));
    InMux I__2317 (
            .O(N__12819),
            .I(N__12813));
    Span4Mux_h I__2316 (
            .O(N__12816),
            .I(N__12810));
    LocalMux I__2315 (
            .O(N__12813),
            .I(N__12807));
    Odrv4 I__2314 (
            .O(N__12810),
            .I(\Lab_UT.sccEldByte ));
    Odrv12 I__2313 (
            .O(N__12807),
            .I(\Lab_UT.sccEldByte ));
    InMux I__2312 (
            .O(N__12802),
            .I(N__12769));
    InMux I__2311 (
            .O(N__12801),
            .I(N__12769));
    InMux I__2310 (
            .O(N__12800),
            .I(N__12769));
    InMux I__2309 (
            .O(N__12799),
            .I(N__12769));
    InMux I__2308 (
            .O(N__12798),
            .I(N__12769));
    InMux I__2307 (
            .O(N__12797),
            .I(N__12769));
    InMux I__2306 (
            .O(N__12796),
            .I(N__12769));
    InMux I__2305 (
            .O(N__12795),
            .I(N__12769));
    InMux I__2304 (
            .O(N__12794),
            .I(N__12752));
    InMux I__2303 (
            .O(N__12793),
            .I(N__12752));
    InMux I__2302 (
            .O(N__12792),
            .I(N__12752));
    InMux I__2301 (
            .O(N__12791),
            .I(N__12752));
    InMux I__2300 (
            .O(N__12790),
            .I(N__12752));
    InMux I__2299 (
            .O(N__12789),
            .I(N__12752));
    InMux I__2298 (
            .O(N__12788),
            .I(N__12752));
    InMux I__2297 (
            .O(N__12787),
            .I(N__12752));
    InMux I__2296 (
            .O(N__12786),
            .I(N__12733));
    LocalMux I__2295 (
            .O(N__12769),
            .I(N__12728));
    LocalMux I__2294 (
            .O(N__12752),
            .I(N__12728));
    InMux I__2293 (
            .O(N__12751),
            .I(N__12713));
    InMux I__2292 (
            .O(N__12750),
            .I(N__12713));
    InMux I__2291 (
            .O(N__12749),
            .I(N__12713));
    InMux I__2290 (
            .O(N__12748),
            .I(N__12713));
    InMux I__2289 (
            .O(N__12747),
            .I(N__12713));
    InMux I__2288 (
            .O(N__12746),
            .I(N__12713));
    InMux I__2287 (
            .O(N__12745),
            .I(N__12713));
    InMux I__2286 (
            .O(N__12744),
            .I(N__12710));
    InMux I__2285 (
            .O(N__12743),
            .I(N__12693));
    InMux I__2284 (
            .O(N__12742),
            .I(N__12693));
    InMux I__2283 (
            .O(N__12741),
            .I(N__12693));
    InMux I__2282 (
            .O(N__12740),
            .I(N__12693));
    InMux I__2281 (
            .O(N__12739),
            .I(N__12693));
    InMux I__2280 (
            .O(N__12738),
            .I(N__12693));
    InMux I__2279 (
            .O(N__12737),
            .I(N__12693));
    InMux I__2278 (
            .O(N__12736),
            .I(N__12693));
    LocalMux I__2277 (
            .O(N__12733),
            .I(N__12688));
    Span4Mux_v I__2276 (
            .O(N__12728),
            .I(N__12688));
    LocalMux I__2275 (
            .O(N__12713),
            .I(N__12683));
    LocalMux I__2274 (
            .O(N__12710),
            .I(N__12683));
    LocalMux I__2273 (
            .O(N__12693),
            .I(\Lab_UT.state_ret_6_RNIL97G01_0 ));
    Odrv4 I__2272 (
            .O(N__12688),
            .I(\Lab_UT.state_ret_6_RNIL97G01_0 ));
    Odrv12 I__2271 (
            .O(N__12683),
            .I(\Lab_UT.state_ret_6_RNIL97G01_0 ));
    IoInMux I__2270 (
            .O(N__12676),
            .I(N__12673));
    LocalMux I__2269 (
            .O(N__12673),
            .I(\Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_iZ0 ));
    CascadeMux I__2268 (
            .O(N__12670),
            .I(\Lab_UT.scctrl.un1_state_inv_cascade_ ));
    CascadeMux I__2267 (
            .O(N__12667),
            .I(\Lab_UT.scctrl.state_ret_12_RNIUQFKZ0_cascade_ ));
    CascadeMux I__2266 (
            .O(N__12664),
            .I(\Lab_UT.state_ret_12_RNIMJCP8_0_cascade_ ));
    InMux I__2265 (
            .O(N__12661),
            .I(N__12658));
    LocalMux I__2264 (
            .O(N__12658),
            .I(\Lab_UT.scctrl.delayload ));
    InMux I__2263 (
            .O(N__12655),
            .I(N__12651));
    InMux I__2262 (
            .O(N__12654),
            .I(N__12648));
    LocalMux I__2261 (
            .O(N__12651),
            .I(N__12645));
    LocalMux I__2260 (
            .O(N__12648),
            .I(N__12640));
    Span4Mux_h I__2259 (
            .O(N__12645),
            .I(N__12640));
    Span4Mux_v I__2258 (
            .O(N__12640),
            .I(N__12637));
    Odrv4 I__2257 (
            .O(N__12637),
            .I(\Lab_UT.scctrl.delay3 ));
    InMux I__2256 (
            .O(N__12634),
            .I(N__12631));
    LocalMux I__2255 (
            .O(N__12631),
            .I(N__12628));
    Odrv4 I__2254 (
            .O(N__12628),
            .I(\Lab_UT.scctrl.r4.delay4 ));
    InMux I__2253 (
            .O(N__12625),
            .I(N__12622));
    LocalMux I__2252 (
            .O(N__12622),
            .I(N__12619));
    Span4Mux_v I__2251 (
            .O(N__12619),
            .I(N__12616));
    Odrv4 I__2250 (
            .O(N__12616),
            .I(\Lab_UT.scdp.u1.byteToDecrypt_2 ));
    InMux I__2249 (
            .O(N__12613),
            .I(N__12609));
    InMux I__2248 (
            .O(N__12612),
            .I(N__12606));
    LocalMux I__2247 (
            .O(N__12609),
            .I(N__12603));
    LocalMux I__2246 (
            .O(N__12606),
            .I(\Lab_UT.scdp.key1_5 ));
    Odrv12 I__2245 (
            .O(N__12603),
            .I(\Lab_UT.scdp.key1_5 ));
    InMux I__2244 (
            .O(N__12598),
            .I(N__12594));
    CascadeMux I__2243 (
            .O(N__12597),
            .I(N__12591));
    LocalMux I__2242 (
            .O(N__12594),
            .I(N__12588));
    InMux I__2241 (
            .O(N__12591),
            .I(N__12585));
    Span4Mux_h I__2240 (
            .O(N__12588),
            .I(N__12582));
    LocalMux I__2239 (
            .O(N__12585),
            .I(\Lab_UT.scdp.key1_1 ));
    Odrv4 I__2238 (
            .O(N__12582),
            .I(\Lab_UT.scdp.key1_1 ));
    InMux I__2237 (
            .O(N__12577),
            .I(N__12574));
    LocalMux I__2236 (
            .O(N__12574),
            .I(N__12570));
    InMux I__2235 (
            .O(N__12573),
            .I(N__12567));
    Span12Mux_s5_h I__2234 (
            .O(N__12570),
            .I(N__12564));
    LocalMux I__2233 (
            .O(N__12567),
            .I(\Lab_UT.scdp.key2_5 ));
    Odrv12 I__2232 (
            .O(N__12564),
            .I(\Lab_UT.scdp.key2_5 ));
    InMux I__2231 (
            .O(N__12559),
            .I(N__12555));
    InMux I__2230 (
            .O(N__12558),
            .I(N__12552));
    LocalMux I__2229 (
            .O(N__12555),
            .I(N__12549));
    LocalMux I__2228 (
            .O(N__12552),
            .I(\Lab_UT.scdp.key3_5 ));
    Odrv4 I__2227 (
            .O(N__12549),
            .I(\Lab_UT.scdp.key3_5 ));
    InMux I__2226 (
            .O(N__12544),
            .I(N__12541));
    LocalMux I__2225 (
            .O(N__12541),
            .I(N__12537));
    InMux I__2224 (
            .O(N__12540),
            .I(N__12534));
    Span4Mux_h I__2223 (
            .O(N__12537),
            .I(N__12531));
    LocalMux I__2222 (
            .O(N__12534),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0 ));
    Odrv4 I__2221 (
            .O(N__12531),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0 ));
    InMux I__2220 (
            .O(N__12526),
            .I(N__12523));
    LocalMux I__2219 (
            .O(N__12523),
            .I(N__12519));
    InMux I__2218 (
            .O(N__12522),
            .I(N__12516));
    Span4Mux_h I__2217 (
            .O(N__12519),
            .I(N__12513));
    LocalMux I__2216 (
            .O(N__12516),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1 ));
    Odrv4 I__2215 (
            .O(N__12513),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1 ));
    InMux I__2214 (
            .O(N__12508),
            .I(N__12504));
    CascadeMux I__2213 (
            .O(N__12507),
            .I(N__12501));
    LocalMux I__2212 (
            .O(N__12504),
            .I(N__12497));
    InMux I__2211 (
            .O(N__12501),
            .I(N__12492));
    InMux I__2210 (
            .O(N__12500),
            .I(N__12492));
    Span4Mux_h I__2209 (
            .O(N__12497),
            .I(N__12489));
    LocalMux I__2208 (
            .O(N__12492),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_12 ));
    Odrv4 I__2207 (
            .O(N__12489),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_12 ));
    InMux I__2206 (
            .O(N__12484),
            .I(N__12480));
    InMux I__2205 (
            .O(N__12483),
            .I(N__12477));
    LocalMux I__2204 (
            .O(N__12480),
            .I(N__12474));
    LocalMux I__2203 (
            .O(N__12477),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13 ));
    Odrv4 I__2202 (
            .O(N__12474),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13 ));
    CEMux I__2201 (
            .O(N__12469),
            .I(N__12457));
    CEMux I__2200 (
            .O(N__12468),
            .I(N__12457));
    CEMux I__2199 (
            .O(N__12467),
            .I(N__12457));
    CEMux I__2198 (
            .O(N__12466),
            .I(N__12457));
    GlobalMux I__2197 (
            .O(N__12457),
            .I(N__12454));
    gio2CtrlBuf I__2196 (
            .O(N__12454),
            .I(\Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_g ));
    InMux I__2195 (
            .O(N__12451),
            .I(N__12447));
    InMux I__2194 (
            .O(N__12450),
            .I(N__12444));
    LocalMux I__2193 (
            .O(N__12447),
            .I(\Lab_UT.scdp.key3_0 ));
    LocalMux I__2192 (
            .O(N__12444),
            .I(\Lab_UT.scdp.key3_0 ));
    InMux I__2191 (
            .O(N__12439),
            .I(N__12436));
    LocalMux I__2190 (
            .O(N__12436),
            .I(N__12431));
    InMux I__2189 (
            .O(N__12435),
            .I(N__12427));
    CascadeMux I__2188 (
            .O(N__12434),
            .I(N__12420));
    Span4Mux_v I__2187 (
            .O(N__12431),
            .I(N__12416));
    InMux I__2186 (
            .O(N__12430),
            .I(N__12413));
    LocalMux I__2185 (
            .O(N__12427),
            .I(N__12410));
    InMux I__2184 (
            .O(N__12426),
            .I(N__12405));
    InMux I__2183 (
            .O(N__12425),
            .I(N__12405));
    InMux I__2182 (
            .O(N__12424),
            .I(N__12400));
    InMux I__2181 (
            .O(N__12423),
            .I(N__12400));
    InMux I__2180 (
            .O(N__12420),
            .I(N__12397));
    InMux I__2179 (
            .O(N__12419),
            .I(N__12394));
    Odrv4 I__2178 (
            .O(N__12416),
            .I(buart__rx_bitcount_2));
    LocalMux I__2177 (
            .O(N__12413),
            .I(buart__rx_bitcount_2));
    Odrv4 I__2176 (
            .O(N__12410),
            .I(buart__rx_bitcount_2));
    LocalMux I__2175 (
            .O(N__12405),
            .I(buart__rx_bitcount_2));
    LocalMux I__2174 (
            .O(N__12400),
            .I(buart__rx_bitcount_2));
    LocalMux I__2173 (
            .O(N__12397),
            .I(buart__rx_bitcount_2));
    LocalMux I__2172 (
            .O(N__12394),
            .I(buart__rx_bitcount_2));
    InMux I__2171 (
            .O(N__12379),
            .I(N__12376));
    LocalMux I__2170 (
            .O(N__12376),
            .I(N__12373));
    Span4Mux_v I__2169 (
            .O(N__12373),
            .I(N__12369));
    InMux I__2168 (
            .O(N__12372),
            .I(N__12366));
    Odrv4 I__2167 (
            .O(N__12369),
            .I(\buart.Z_rx.bitcount_es_RNIGTPI1Z0Z_3 ));
    LocalMux I__2166 (
            .O(N__12366),
            .I(\buart.Z_rx.bitcount_es_RNIGTPI1Z0Z_3 ));
    InMux I__2165 (
            .O(N__12361),
            .I(N__12358));
    LocalMux I__2164 (
            .O(N__12358),
            .I(N__12353));
    InMux I__2163 (
            .O(N__12357),
            .I(N__12348));
    InMux I__2162 (
            .O(N__12356),
            .I(N__12348));
    Span4Mux_h I__2161 (
            .O(N__12353),
            .I(N__12345));
    LocalMux I__2160 (
            .O(N__12348),
            .I(N__12342));
    Odrv4 I__2159 (
            .O(N__12345),
            .I(\Lab_UT.scdp.d2eData_0 ));
    Odrv4 I__2158 (
            .O(N__12342),
            .I(\Lab_UT.scdp.d2eData_0 ));
    InMux I__2157 (
            .O(N__12337),
            .I(N__12334));
    LocalMux I__2156 (
            .O(N__12334),
            .I(N__12330));
    CascadeMux I__2155 (
            .O(N__12333),
            .I(N__12327));
    Span4Mux_v I__2154 (
            .O(N__12330),
            .I(N__12324));
    InMux I__2153 (
            .O(N__12327),
            .I(N__12321));
    Span4Mux_v I__2152 (
            .O(N__12324),
            .I(N__12318));
    LocalMux I__2151 (
            .O(N__12321),
            .I(\Lab_UT.scdp.lsBitsD_0 ));
    Odrv4 I__2150 (
            .O(N__12318),
            .I(\Lab_UT.scdp.lsBitsD_0 ));
    InMux I__2149 (
            .O(N__12313),
            .I(N__12309));
    InMux I__2148 (
            .O(N__12312),
            .I(N__12306));
    LocalMux I__2147 (
            .O(N__12309),
            .I(N__12299));
    LocalMux I__2146 (
            .O(N__12306),
            .I(N__12299));
    InMux I__2145 (
            .O(N__12305),
            .I(N__12294));
    InMux I__2144 (
            .O(N__12304),
            .I(N__12294));
    Span4Mux_h I__2143 (
            .O(N__12299),
            .I(N__12291));
    LocalMux I__2142 (
            .O(N__12294),
            .I(\Lab_UT.scdp.lsBits_6 ));
    Odrv4 I__2141 (
            .O(N__12291),
            .I(\Lab_UT.scdp.lsBits_6 ));
    InMux I__2140 (
            .O(N__12286),
            .I(N__12282));
    InMux I__2139 (
            .O(N__12285),
            .I(N__12279));
    LocalMux I__2138 (
            .O(N__12282),
            .I(N__12276));
    LocalMux I__2137 (
            .O(N__12279),
            .I(N__12271));
    Span4Mux_s3_v I__2136 (
            .O(N__12276),
            .I(N__12271));
    Odrv4 I__2135 (
            .O(N__12271),
            .I(\Lab_UT.scdp.lsBitsD_4 ));
    InMux I__2134 (
            .O(N__12268),
            .I(N__12264));
    CascadeMux I__2133 (
            .O(N__12267),
            .I(N__12260));
    LocalMux I__2132 (
            .O(N__12264),
            .I(N__12255));
    InMux I__2131 (
            .O(N__12263),
            .I(N__12248));
    InMux I__2130 (
            .O(N__12260),
            .I(N__12248));
    InMux I__2129 (
            .O(N__12259),
            .I(N__12248));
    InMux I__2128 (
            .O(N__12258),
            .I(N__12245));
    Span4Mux_h I__2127 (
            .O(N__12255),
            .I(N__12242));
    LocalMux I__2126 (
            .O(N__12248),
            .I(N__12237));
    LocalMux I__2125 (
            .O(N__12245),
            .I(N__12237));
    Span4Mux_v I__2124 (
            .O(N__12242),
            .I(N__12232));
    Span4Mux_v I__2123 (
            .O(N__12237),
            .I(N__12232));
    Odrv4 I__2122 (
            .O(N__12232),
            .I(\Lab_UT.scdp.N_48_i ));
    InMux I__2121 (
            .O(N__12229),
            .I(N__12226));
    LocalMux I__2120 (
            .O(N__12226),
            .I(N__12223));
    Span4Mux_v I__2119 (
            .O(N__12223),
            .I(N__12220));
    Span4Mux_v I__2118 (
            .O(N__12220),
            .I(N__12216));
    InMux I__2117 (
            .O(N__12219),
            .I(N__12213));
    Odrv4 I__2116 (
            .O(N__12216),
            .I(\Lab_UT.scdp.N_52 ));
    LocalMux I__2115 (
            .O(N__12213),
            .I(\Lab_UT.scdp.N_52 ));
    InMux I__2114 (
            .O(N__12208),
            .I(N__12204));
    CascadeMux I__2113 (
            .O(N__12207),
            .I(N__12201));
    LocalMux I__2112 (
            .O(N__12204),
            .I(N__12198));
    InMux I__2111 (
            .O(N__12201),
            .I(N__12195));
    Span4Mux_h I__2110 (
            .O(N__12198),
            .I(N__12192));
    LocalMux I__2109 (
            .O(N__12195),
            .I(N__12187));
    Span4Mux_v I__2108 (
            .O(N__12192),
            .I(N__12187));
    Odrv4 I__2107 (
            .O(N__12187),
            .I(\Lab_UT.scdp.msBitsD_3 ));
    InMux I__2106 (
            .O(N__12184),
            .I(N__12181));
    LocalMux I__2105 (
            .O(N__12181),
            .I(N__12172));
    InMux I__2104 (
            .O(N__12180),
            .I(N__12169));
    InMux I__2103 (
            .O(N__12179),
            .I(N__12166));
    InMux I__2102 (
            .O(N__12178),
            .I(N__12159));
    InMux I__2101 (
            .O(N__12177),
            .I(N__12159));
    InMux I__2100 (
            .O(N__12176),
            .I(N__12159));
    InMux I__2099 (
            .O(N__12175),
            .I(N__12155));
    Span4Mux_h I__2098 (
            .O(N__12172),
            .I(N__12152));
    LocalMux I__2097 (
            .O(N__12169),
            .I(N__12149));
    LocalMux I__2096 (
            .O(N__12166),
            .I(N__12146));
    LocalMux I__2095 (
            .O(N__12159),
            .I(N__12143));
    InMux I__2094 (
            .O(N__12158),
            .I(N__12140));
    LocalMux I__2093 (
            .O(N__12155),
            .I(N__12137));
    Span4Mux_v I__2092 (
            .O(N__12152),
            .I(N__12132));
    Span4Mux_h I__2091 (
            .O(N__12149),
            .I(N__12132));
    Span4Mux_v I__2090 (
            .O(N__12146),
            .I(N__12127));
    Span4Mux_v I__2089 (
            .O(N__12143),
            .I(N__12127));
    LocalMux I__2088 (
            .O(N__12140),
            .I(N__12124));
    Odrv4 I__2087 (
            .O(N__12137),
            .I(buart__tx_uart_busy_0_i));
    Odrv4 I__2086 (
            .O(N__12132),
            .I(buart__tx_uart_busy_0_i));
    Odrv4 I__2085 (
            .O(N__12127),
            .I(buart__tx_uart_busy_0_i));
    Odrv4 I__2084 (
            .O(N__12124),
            .I(buart__tx_uart_busy_0_i));
    CascadeMux I__2083 (
            .O(N__12115),
            .I(N__12112));
    InMux I__2082 (
            .O(N__12112),
            .I(N__12109));
    LocalMux I__2081 (
            .O(N__12109),
            .I(N__12106));
    Span4Mux_v I__2080 (
            .O(N__12106),
            .I(N__12100));
    InMux I__2079 (
            .O(N__12105),
            .I(N__12097));
    CascadeMux I__2078 (
            .O(N__12104),
            .I(N__12090));
    CascadeMux I__2077 (
            .O(N__12103),
            .I(N__12087));
    Span4Mux_h I__2076 (
            .O(N__12100),
            .I(N__12081));
    LocalMux I__2075 (
            .O(N__12097),
            .I(N__12081));
    InMux I__2074 (
            .O(N__12096),
            .I(N__12078));
    InMux I__2073 (
            .O(N__12095),
            .I(N__12071));
    InMux I__2072 (
            .O(N__12094),
            .I(N__12071));
    InMux I__2071 (
            .O(N__12093),
            .I(N__12071));
    InMux I__2070 (
            .O(N__12090),
            .I(N__12064));
    InMux I__2069 (
            .O(N__12087),
            .I(N__12064));
    InMux I__2068 (
            .O(N__12086),
            .I(N__12064));
    Span4Mux_v I__2067 (
            .O(N__12081),
            .I(N__12059));
    LocalMux I__2066 (
            .O(N__12078),
            .I(N__12059));
    LocalMux I__2065 (
            .O(N__12071),
            .I(\buart.Z_tx.N_255 ));
    LocalMux I__2064 (
            .O(N__12064),
            .I(\buart.Z_tx.N_255 ));
    Odrv4 I__2063 (
            .O(N__12059),
            .I(\buart.Z_tx.N_255 ));
    InMux I__2062 (
            .O(N__12052),
            .I(N__12044));
    InMux I__2061 (
            .O(N__12051),
            .I(N__12030));
    InMux I__2060 (
            .O(N__12050),
            .I(N__12030));
    InMux I__2059 (
            .O(N__12049),
            .I(N__12025));
    InMux I__2058 (
            .O(N__12048),
            .I(N__12025));
    InMux I__2057 (
            .O(N__12047),
            .I(N__12022));
    LocalMux I__2056 (
            .O(N__12044),
            .I(N__12019));
    InMux I__2055 (
            .O(N__12043),
            .I(N__12012));
    InMux I__2054 (
            .O(N__12042),
            .I(N__12012));
    InMux I__2053 (
            .O(N__12041),
            .I(N__12012));
    InMux I__2052 (
            .O(N__12040),
            .I(N__12009));
    InMux I__2051 (
            .O(N__12039),
            .I(N__12002));
    InMux I__2050 (
            .O(N__12038),
            .I(N__12002));
    InMux I__2049 (
            .O(N__12037),
            .I(N__12002));
    InMux I__2048 (
            .O(N__12036),
            .I(N__11997));
    InMux I__2047 (
            .O(N__12035),
            .I(N__11997));
    LocalMux I__2046 (
            .O(N__12030),
            .I(N__11994));
    LocalMux I__2045 (
            .O(N__12025),
            .I(N__11989));
    LocalMux I__2044 (
            .O(N__12022),
            .I(N__11989));
    Span12Mux_s9_v I__2043 (
            .O(N__12019),
            .I(N__11986));
    LocalMux I__2042 (
            .O(N__12012),
            .I(N__11981));
    LocalMux I__2041 (
            .O(N__12009),
            .I(N__11981));
    LocalMux I__2040 (
            .O(N__12002),
            .I(ufifo_utb_txdata_rdy_0));
    LocalMux I__2039 (
            .O(N__11997),
            .I(ufifo_utb_txdata_rdy_0));
    Odrv4 I__2038 (
            .O(N__11994),
            .I(ufifo_utb_txdata_rdy_0));
    Odrv4 I__2037 (
            .O(N__11989),
            .I(ufifo_utb_txdata_rdy_0));
    Odrv12 I__2036 (
            .O(N__11986),
            .I(ufifo_utb_txdata_rdy_0));
    Odrv4 I__2035 (
            .O(N__11981),
            .I(ufifo_utb_txdata_rdy_0));
    InMux I__2034 (
            .O(N__11968),
            .I(N__11965));
    LocalMux I__2033 (
            .O(N__11965),
            .I(N__11961));
    InMux I__2032 (
            .O(N__11964),
            .I(N__11957));
    Span4Mux_h I__2031 (
            .O(N__11961),
            .I(N__11954));
    InMux I__2030 (
            .O(N__11960),
            .I(N__11951));
    LocalMux I__2029 (
            .O(N__11957),
            .I(N__11948));
    Span4Mux_v I__2028 (
            .O(N__11954),
            .I(N__11945));
    LocalMux I__2027 (
            .O(N__11951),
            .I(N__11940));
    Span12Mux_v I__2026 (
            .O(N__11948),
            .I(N__11940));
    Odrv4 I__2025 (
            .O(N__11945),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    Odrv12 I__2024 (
            .O(N__11940),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    CascadeMux I__2023 (
            .O(N__11935),
            .I(N__11929));
    InMux I__2022 (
            .O(N__11934),
            .I(N__11926));
    InMux I__2021 (
            .O(N__11933),
            .I(N__11914));
    InMux I__2020 (
            .O(N__11932),
            .I(N__11914));
    InMux I__2019 (
            .O(N__11929),
            .I(N__11914));
    LocalMux I__2018 (
            .O(N__11926),
            .I(N__11911));
    InMux I__2017 (
            .O(N__11925),
            .I(N__11904));
    InMux I__2016 (
            .O(N__11924),
            .I(N__11904));
    InMux I__2015 (
            .O(N__11923),
            .I(N__11904));
    InMux I__2014 (
            .O(N__11922),
            .I(N__11899));
    InMux I__2013 (
            .O(N__11921),
            .I(N__11899));
    LocalMux I__2012 (
            .O(N__11914),
            .I(N__11894));
    Span4Mux_v I__2011 (
            .O(N__11911),
            .I(N__11887));
    LocalMux I__2010 (
            .O(N__11904),
            .I(N__11887));
    LocalMux I__2009 (
            .O(N__11899),
            .I(N__11887));
    InMux I__2008 (
            .O(N__11898),
            .I(N__11882));
    InMux I__2007 (
            .O(N__11897),
            .I(N__11882));
    Span4Mux_v I__2006 (
            .O(N__11894),
            .I(N__11877));
    Span4Mux_h I__2005 (
            .O(N__11887),
            .I(N__11877));
    LocalMux I__2004 (
            .O(N__11882),
            .I(bu_rx_data_3));
    Odrv4 I__2003 (
            .O(N__11877),
            .I(bu_rx_data_3));
    CascadeMux I__2002 (
            .O(N__11872),
            .I(\Lab_UT.scdp.a2b.N_53_cascade_ ));
    InMux I__2001 (
            .O(N__11869),
            .I(N__11866));
    LocalMux I__2000 (
            .O(N__11866),
            .I(N__11862));
    InMux I__1999 (
            .O(N__11865),
            .I(N__11859));
    Span4Mux_h I__1998 (
            .O(N__11862),
            .I(N__11856));
    LocalMux I__1997 (
            .O(N__11859),
            .I(N__11851));
    Span4Mux_v I__1996 (
            .O(N__11856),
            .I(N__11851));
    Odrv4 I__1995 (
            .O(N__11851),
            .I(\Lab_UT.scdp.N_39 ));
    CascadeMux I__1994 (
            .O(N__11848),
            .I(N__11844));
    InMux I__1993 (
            .O(N__11847),
            .I(N__11839));
    InMux I__1992 (
            .O(N__11844),
            .I(N__11839));
    LocalMux I__1991 (
            .O(N__11839),
            .I(N__11835));
    InMux I__1990 (
            .O(N__11838),
            .I(N__11832));
    Span4Mux_h I__1989 (
            .O(N__11835),
            .I(N__11829));
    LocalMux I__1988 (
            .O(N__11832),
            .I(\Lab_UT.scdp.byteToDecrypt_4 ));
    Odrv4 I__1987 (
            .O(N__11829),
            .I(\Lab_UT.scdp.byteToDecrypt_4 ));
    InMux I__1986 (
            .O(N__11824),
            .I(N__11820));
    CascadeMux I__1985 (
            .O(N__11823),
            .I(N__11816));
    LocalMux I__1984 (
            .O(N__11820),
            .I(N__11813));
    InMux I__1983 (
            .O(N__11819),
            .I(N__11810));
    InMux I__1982 (
            .O(N__11816),
            .I(N__11807));
    Span4Mux_h I__1981 (
            .O(N__11813),
            .I(N__11804));
    LocalMux I__1980 (
            .O(N__11810),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_6 ));
    LocalMux I__1979 (
            .O(N__11807),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_6 ));
    Odrv4 I__1978 (
            .O(N__11804),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_6 ));
    CascadeMux I__1977 (
            .O(N__11797),
            .I(N__11793));
    InMux I__1976 (
            .O(N__11796),
            .I(N__11790));
    InMux I__1975 (
            .O(N__11793),
            .I(N__11787));
    LocalMux I__1974 (
            .O(N__11790),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30 ));
    LocalMux I__1973 (
            .O(N__11787),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30 ));
    CascadeMux I__1972 (
            .O(N__11782),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsr_next_1_0_cascade_ ));
    InMux I__1971 (
            .O(N__11779),
            .I(N__11774));
    InMux I__1970 (
            .O(N__11778),
            .I(N__11771));
    InMux I__1969 (
            .O(N__11777),
            .I(N__11768));
    LocalMux I__1968 (
            .O(N__11774),
            .I(N__11765));
    LocalMux I__1967 (
            .O(N__11771),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2 ));
    LocalMux I__1966 (
            .O(N__11768),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2 ));
    Odrv4 I__1965 (
            .O(N__11765),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2 ));
    InMux I__1964 (
            .O(N__11758),
            .I(N__11754));
    InMux I__1963 (
            .O(N__11757),
            .I(N__11751));
    LocalMux I__1962 (
            .O(N__11754),
            .I(N__11748));
    LocalMux I__1961 (
            .O(N__11751),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_4 ));
    Odrv4 I__1960 (
            .O(N__11748),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_4 ));
    InMux I__1959 (
            .O(N__11743),
            .I(N__11738));
    InMux I__1958 (
            .O(N__11742),
            .I(N__11733));
    InMux I__1957 (
            .O(N__11741),
            .I(N__11733));
    LocalMux I__1956 (
            .O(N__11738),
            .I(N__11730));
    LocalMux I__1955 (
            .O(N__11733),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5 ));
    Odrv4 I__1954 (
            .O(N__11730),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5 ));
    InMux I__1953 (
            .O(N__11725),
            .I(N__11721));
    InMux I__1952 (
            .O(N__11724),
            .I(N__11718));
    LocalMux I__1951 (
            .O(N__11721),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_11 ));
    LocalMux I__1950 (
            .O(N__11718),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_11 ));
    InMux I__1949 (
            .O(N__11713),
            .I(N__11710));
    LocalMux I__1948 (
            .O(N__11710),
            .I(\Lab_UT.scctrl.next_state_0_sqmuxa_4Z0Z_0 ));
    InMux I__1947 (
            .O(N__11707),
            .I(N__11704));
    LocalMux I__1946 (
            .O(N__11704),
            .I(\Lab_UT.dk.de_bigEZ0Z_1 ));
    CascadeMux I__1945 (
            .O(N__11701),
            .I(Lab_UT_dk_de_bigD_6_cascade_));
    CascadeMux I__1944 (
            .O(N__11698),
            .I(\Lab_UT.de_bigE_cascade_ ));
    CascadeMux I__1943 (
            .O(N__11695),
            .I(\Lab_UT.scdp.N_39_cascade_ ));
    CascadeMux I__1942 (
            .O(N__11692),
            .I(\Lab_UT.scdp.a2b.N_50_cascade_ ));
    CascadeMux I__1941 (
            .O(N__11689),
            .I(N__11686));
    InMux I__1940 (
            .O(N__11686),
            .I(N__11683));
    LocalMux I__1939 (
            .O(N__11683),
            .I(\Lab_UT.scdp.a2b.N_51 ));
    InMux I__1938 (
            .O(N__11680),
            .I(N__11675));
    InMux I__1937 (
            .O(N__11679),
            .I(N__11669));
    InMux I__1936 (
            .O(N__11678),
            .I(N__11669));
    LocalMux I__1935 (
            .O(N__11675),
            .I(N__11666));
    CascadeMux I__1934 (
            .O(N__11674),
            .I(N__11662));
    LocalMux I__1933 (
            .O(N__11669),
            .I(N__11659));
    Span4Mux_h I__1932 (
            .O(N__11666),
            .I(N__11656));
    InMux I__1931 (
            .O(N__11665),
            .I(N__11653));
    InMux I__1930 (
            .O(N__11662),
            .I(N__11650));
    Odrv4 I__1929 (
            .O(N__11659),
            .I(bu_rx_data_i_2_5));
    Odrv4 I__1928 (
            .O(N__11656),
            .I(bu_rx_data_i_2_5));
    LocalMux I__1927 (
            .O(N__11653),
            .I(bu_rx_data_i_2_5));
    LocalMux I__1926 (
            .O(N__11650),
            .I(bu_rx_data_i_2_5));
    CascadeMux I__1925 (
            .O(N__11641),
            .I(N__11638));
    InMux I__1924 (
            .O(N__11638),
            .I(N__11635));
    LocalMux I__1923 (
            .O(N__11635),
            .I(N__11632));
    Span4Mux_h I__1922 (
            .O(N__11632),
            .I(N__11629));
    Odrv4 I__1921 (
            .O(N__11629),
            .I(\Lab_UT.scctrl.m24_e_5 ));
    InMux I__1920 (
            .O(N__11626),
            .I(N__11623));
    LocalMux I__1919 (
            .O(N__11623),
            .I(N__11620));
    Span4Mux_v I__1918 (
            .O(N__11620),
            .I(N__11616));
    InMux I__1917 (
            .O(N__11619),
            .I(N__11613));
    Odrv4 I__1916 (
            .O(N__11616),
            .I(\Lab_UT.scdp.a2b.N_50 ));
    LocalMux I__1915 (
            .O(N__11613),
            .I(\Lab_UT.scdp.a2b.N_50 ));
    CascadeMux I__1914 (
            .O(N__11608),
            .I(bu_rx_data_rdy_cascade_));
    InMux I__1913 (
            .O(N__11605),
            .I(N__11602));
    LocalMux I__1912 (
            .O(N__11602),
            .I(\Lab_UT.scctrl.delay1 ));
    InMux I__1911 (
            .O(N__11599),
            .I(N__11596));
    LocalMux I__1910 (
            .O(N__11596),
            .I(\Lab_UT.scctrl.delay2 ));
    InMux I__1909 (
            .O(N__11593),
            .I(N__11587));
    InMux I__1908 (
            .O(N__11592),
            .I(N__11587));
    LocalMux I__1907 (
            .O(N__11587),
            .I(N__11583));
    InMux I__1906 (
            .O(N__11586),
            .I(N__11580));
    Span4Mux_v I__1905 (
            .O(N__11583),
            .I(N__11575));
    LocalMux I__1904 (
            .O(N__11580),
            .I(N__11575));
    Odrv4 I__1903 (
            .O(N__11575),
            .I(N_6));
    CascadeMux I__1902 (
            .O(N__11572),
            .I(\Lab_UT.scdp.pinst1.un12_pValidZ0Z_1_cascade_ ));
    InMux I__1901 (
            .O(N__11569),
            .I(N__11566));
    LocalMux I__1900 (
            .O(N__11566),
            .I(\Lab_UT.un7_pValid ));
    InMux I__1899 (
            .O(N__11563),
            .I(N__11557));
    InMux I__1898 (
            .O(N__11562),
            .I(N__11557));
    LocalMux I__1897 (
            .O(N__11557),
            .I(\Lab_UT.un1_pValid ));
    CascadeMux I__1896 (
            .O(N__11554),
            .I(\Lab_UT.un7_pValid_cascade_ ));
    CascadeMux I__1895 (
            .O(N__11551),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_1_0_i_cascade_ ));
    CascadeMux I__1894 (
            .O(N__11548),
            .I(\Lab_UT.g0_i_a9_1_3_cascade_ ));
    InMux I__1893 (
            .O(N__11545),
            .I(N__11542));
    LocalMux I__1892 (
            .O(N__11542),
            .I(\Lab_UT.scctrl.m24_e_4 ));
    CascadeMux I__1891 (
            .O(N__11539),
            .I(\Lab_UT.dk.escKey_4_reti_cascade_ ));
    InMux I__1890 (
            .O(N__11536),
            .I(N__11533));
    LocalMux I__1889 (
            .O(N__11533),
            .I(N__11530));
    Odrv4 I__1888 (
            .O(N__11530),
            .I(\Lab_UT.scctrl.g0_i_a7_1 ));
    CascadeMux I__1887 (
            .O(N__11527),
            .I(\Lab_UT.scctrl.g0_i_a3_2_cascade_ ));
    InMux I__1886 (
            .O(N__11524),
            .I(N__11520));
    CascadeMux I__1885 (
            .O(N__11523),
            .I(N__11514));
    LocalMux I__1884 (
            .O(N__11520),
            .I(N__11510));
    InMux I__1883 (
            .O(N__11519),
            .I(N__11507));
    InMux I__1882 (
            .O(N__11518),
            .I(N__11504));
    InMux I__1881 (
            .O(N__11517),
            .I(N__11501));
    InMux I__1880 (
            .O(N__11514),
            .I(N__11496));
    InMux I__1879 (
            .O(N__11513),
            .I(N__11496));
    Odrv4 I__1878 (
            .O(N__11510),
            .I(\ufifo.tx_fsm.cstateZ0Z_4 ));
    LocalMux I__1877 (
            .O(N__11507),
            .I(\ufifo.tx_fsm.cstateZ0Z_4 ));
    LocalMux I__1876 (
            .O(N__11504),
            .I(\ufifo.tx_fsm.cstateZ0Z_4 ));
    LocalMux I__1875 (
            .O(N__11501),
            .I(\ufifo.tx_fsm.cstateZ0Z_4 ));
    LocalMux I__1874 (
            .O(N__11496),
            .I(\ufifo.tx_fsm.cstateZ0Z_4 ));
    InMux I__1873 (
            .O(N__11485),
            .I(N__11481));
    InMux I__1872 (
            .O(N__11484),
            .I(N__11478));
    LocalMux I__1871 (
            .O(N__11481),
            .I(\ufifo.tx_fsm.N_59_0 ));
    LocalMux I__1870 (
            .O(N__11478),
            .I(\ufifo.tx_fsm.N_59_0 ));
    InMux I__1869 (
            .O(N__11473),
            .I(N__11470));
    LocalMux I__1868 (
            .O(N__11470),
            .I(N__11464));
    InMux I__1867 (
            .O(N__11469),
            .I(N__11459));
    InMux I__1866 (
            .O(N__11468),
            .I(N__11456));
    InMux I__1865 (
            .O(N__11467),
            .I(N__11453));
    Span4Mux_v I__1864 (
            .O(N__11464),
            .I(N__11449));
    InMux I__1863 (
            .O(N__11463),
            .I(N__11444));
    InMux I__1862 (
            .O(N__11462),
            .I(N__11444));
    LocalMux I__1861 (
            .O(N__11459),
            .I(N__11439));
    LocalMux I__1860 (
            .O(N__11456),
            .I(N__11436));
    LocalMux I__1859 (
            .O(N__11453),
            .I(N__11433));
    InMux I__1858 (
            .O(N__11452),
            .I(N__11429));
    Sp12to4 I__1857 (
            .O(N__11449),
            .I(N__11424));
    LocalMux I__1856 (
            .O(N__11444),
            .I(N__11424));
    InMux I__1855 (
            .O(N__11443),
            .I(N__11419));
    InMux I__1854 (
            .O(N__11442),
            .I(N__11419));
    Span4Mux_h I__1853 (
            .O(N__11439),
            .I(N__11416));
    Span4Mux_v I__1852 (
            .O(N__11436),
            .I(N__11411));
    Span4Mux_h I__1851 (
            .O(N__11433),
            .I(N__11411));
    InMux I__1850 (
            .O(N__11432),
            .I(N__11408));
    LocalMux I__1849 (
            .O(N__11429),
            .I(buart__tx_uart_busy_0));
    Odrv12 I__1848 (
            .O(N__11424),
            .I(buart__tx_uart_busy_0));
    LocalMux I__1847 (
            .O(N__11419),
            .I(buart__tx_uart_busy_0));
    Odrv4 I__1846 (
            .O(N__11416),
            .I(buart__tx_uart_busy_0));
    Odrv4 I__1845 (
            .O(N__11411),
            .I(buart__tx_uart_busy_0));
    LocalMux I__1844 (
            .O(N__11408),
            .I(buart__tx_uart_busy_0));
    InMux I__1843 (
            .O(N__11395),
            .I(N__11391));
    InMux I__1842 (
            .O(N__11394),
            .I(N__11388));
    LocalMux I__1841 (
            .O(N__11391),
            .I(N__11382));
    LocalMux I__1840 (
            .O(N__11388),
            .I(N__11379));
    InMux I__1839 (
            .O(N__11387),
            .I(N__11376));
    InMux I__1838 (
            .O(N__11386),
            .I(N__11371));
    CascadeMux I__1837 (
            .O(N__11385),
            .I(N__11367));
    Span4Mux_h I__1836 (
            .O(N__11382),
            .I(N__11364));
    Span4Mux_v I__1835 (
            .O(N__11379),
            .I(N__11359));
    LocalMux I__1834 (
            .O(N__11376),
            .I(N__11359));
    InMux I__1833 (
            .O(N__11375),
            .I(N__11354));
    InMux I__1832 (
            .O(N__11374),
            .I(N__11354));
    LocalMux I__1831 (
            .O(N__11371),
            .I(N__11351));
    InMux I__1830 (
            .O(N__11370),
            .I(N__11348));
    InMux I__1829 (
            .O(N__11367),
            .I(N__11345));
    Span4Mux_v I__1828 (
            .O(N__11364),
            .I(N__11340));
    Span4Mux_h I__1827 (
            .O(N__11359),
            .I(N__11340));
    LocalMux I__1826 (
            .O(N__11354),
            .I(N__11335));
    Span12Mux_s11_v I__1825 (
            .O(N__11351),
            .I(N__11335));
    LocalMux I__1824 (
            .O(N__11348),
            .I(\ufifo.emitcrlf_fsm.cstateZ0Z_1 ));
    LocalMux I__1823 (
            .O(N__11345),
            .I(\ufifo.emitcrlf_fsm.cstateZ0Z_1 ));
    Odrv4 I__1822 (
            .O(N__11340),
            .I(\ufifo.emitcrlf_fsm.cstateZ0Z_1 ));
    Odrv12 I__1821 (
            .O(N__11335),
            .I(\ufifo.emitcrlf_fsm.cstateZ0Z_1 ));
    InMux I__1820 (
            .O(N__11326),
            .I(N__11323));
    LocalMux I__1819 (
            .O(N__11323),
            .I(\ufifo.emitcrlf_fsm.cstate_srsts_rn_0_1 ));
    InMux I__1818 (
            .O(N__11320),
            .I(N__11316));
    CascadeMux I__1817 (
            .O(N__11319),
            .I(N__11313));
    LocalMux I__1816 (
            .O(N__11316),
            .I(N__11310));
    InMux I__1815 (
            .O(N__11313),
            .I(N__11307));
    Odrv4 I__1814 (
            .O(N__11310),
            .I(\ufifo.tx_fsm.cstateZ0Z_5 ));
    LocalMux I__1813 (
            .O(N__11307),
            .I(\ufifo.tx_fsm.cstateZ0Z_5 ));
    InMux I__1812 (
            .O(N__11302),
            .I(N__11298));
    InMux I__1811 (
            .O(N__11301),
            .I(N__11295));
    LocalMux I__1810 (
            .O(N__11298),
            .I(N__11288));
    LocalMux I__1809 (
            .O(N__11295),
            .I(N__11288));
    InMux I__1808 (
            .O(N__11294),
            .I(N__11283));
    InMux I__1807 (
            .O(N__11293),
            .I(N__11283));
    Span4Mux_v I__1806 (
            .O(N__11288),
            .I(N__11278));
    LocalMux I__1805 (
            .O(N__11283),
            .I(N__11278));
    Span4Mux_h I__1804 (
            .O(N__11278),
            .I(N__11275));
    Odrv4 I__1803 (
            .O(N__11275),
            .I(\ufifo.crlfdone ));
    CascadeMux I__1802 (
            .O(N__11272),
            .I(\ufifo.tx_fsm.N_72_cascade_ ));
    InMux I__1801 (
            .O(N__11269),
            .I(N__11257));
    InMux I__1800 (
            .O(N__11268),
            .I(N__11257));
    InMux I__1799 (
            .O(N__11267),
            .I(N__11246));
    InMux I__1798 (
            .O(N__11266),
            .I(N__11246));
    InMux I__1797 (
            .O(N__11265),
            .I(N__11246));
    InMux I__1796 (
            .O(N__11264),
            .I(N__11246));
    InMux I__1795 (
            .O(N__11263),
            .I(N__11246));
    InMux I__1794 (
            .O(N__11262),
            .I(N__11243));
    LocalMux I__1793 (
            .O(N__11257),
            .I(N__11238));
    LocalMux I__1792 (
            .O(N__11246),
            .I(N__11233));
    LocalMux I__1791 (
            .O(N__11243),
            .I(N__11233));
    InMux I__1790 (
            .O(N__11242),
            .I(N__11230));
    InMux I__1789 (
            .O(N__11241),
            .I(N__11227));
    Span4Mux_v I__1788 (
            .O(N__11238),
            .I(N__11218));
    Span4Mux_v I__1787 (
            .O(N__11233),
            .I(N__11218));
    LocalMux I__1786 (
            .O(N__11230),
            .I(N__11218));
    LocalMux I__1785 (
            .O(N__11227),
            .I(N__11215));
    InMux I__1784 (
            .O(N__11226),
            .I(N__11210));
    InMux I__1783 (
            .O(N__11225),
            .I(N__11210));
    Span4Mux_h I__1782 (
            .O(N__11218),
            .I(N__11207));
    Odrv4 I__1781 (
            .O(N__11215),
            .I(\ufifo.cstate_0 ));
    LocalMux I__1780 (
            .O(N__11210),
            .I(\ufifo.cstate_0 ));
    Odrv4 I__1779 (
            .O(N__11207),
            .I(\ufifo.cstate_0 ));
    InMux I__1778 (
            .O(N__11200),
            .I(N__11197));
    LocalMux I__1777 (
            .O(N__11197),
            .I(\Lab_UT.dk.de_bigEZ0Z_2 ));
    CascadeMux I__1776 (
            .O(N__11194),
            .I(\Lab_UT.scdp.d2eData_3_5_cascade_ ));
    InMux I__1775 (
            .O(N__11191),
            .I(N__11188));
    LocalMux I__1774 (
            .O(N__11188),
            .I(N__11185));
    Span4Mux_h I__1773 (
            .O(N__11185),
            .I(N__11180));
    InMux I__1772 (
            .O(N__11184),
            .I(N__11175));
    InMux I__1771 (
            .O(N__11183),
            .I(N__11175));
    Odrv4 I__1770 (
            .O(N__11180),
            .I(\Lab_UT.scdp.e2dData_5 ));
    LocalMux I__1769 (
            .O(N__11175),
            .I(\Lab_UT.scdp.e2dData_5 ));
    InMux I__1768 (
            .O(N__11170),
            .I(N__11164));
    InMux I__1767 (
            .O(N__11169),
            .I(N__11164));
    LocalMux I__1766 (
            .O(N__11164),
            .I(\Lab_UT.scdp.u0.byteToDecrypt_5 ));
    InMux I__1765 (
            .O(N__11161),
            .I(N__11157));
    InMux I__1764 (
            .O(N__11160),
            .I(N__11154));
    LocalMux I__1763 (
            .O(N__11157),
            .I(\Lab_UT.scdp.u0.byteToDecrypt_7 ));
    LocalMux I__1762 (
            .O(N__11154),
            .I(\Lab_UT.scdp.u0.byteToDecrypt_7 ));
    InMux I__1761 (
            .O(N__11149),
            .I(N__11144));
    InMux I__1760 (
            .O(N__11148),
            .I(N__11141));
    InMux I__1759 (
            .O(N__11147),
            .I(N__11138));
    LocalMux I__1758 (
            .O(N__11144),
            .I(N__11131));
    LocalMux I__1757 (
            .O(N__11141),
            .I(N__11131));
    LocalMux I__1756 (
            .O(N__11138),
            .I(N__11131));
    Span4Mux_v I__1755 (
            .O(N__11131),
            .I(N__11128));
    Odrv4 I__1754 (
            .O(N__11128),
            .I(\Lab_UT.scdp.val_0_3 ));
    InMux I__1753 (
            .O(N__11125),
            .I(N__11122));
    LocalMux I__1752 (
            .O(N__11122),
            .I(N__11118));
    InMux I__1751 (
            .O(N__11121),
            .I(N__11115));
    Span4Mux_h I__1750 (
            .O(N__11118),
            .I(N__11112));
    LocalMux I__1749 (
            .O(N__11115),
            .I(\Lab_UT.scdp.key1_7 ));
    Odrv4 I__1748 (
            .O(N__11112),
            .I(\Lab_UT.scdp.key1_7 ));
    InMux I__1747 (
            .O(N__11107),
            .I(N__11103));
    InMux I__1746 (
            .O(N__11106),
            .I(N__11100));
    LocalMux I__1745 (
            .O(N__11103),
            .I(N__11097));
    LocalMux I__1744 (
            .O(N__11100),
            .I(\Lab_UT.scdp.key1_3 ));
    Odrv12 I__1743 (
            .O(N__11097),
            .I(\Lab_UT.scdp.key1_3 ));
    SRMux I__1742 (
            .O(N__11092),
            .I(N__11087));
    CEMux I__1741 (
            .O(N__11091),
            .I(N__11084));
    CascadeMux I__1740 (
            .O(N__11090),
            .I(N__11080));
    LocalMux I__1739 (
            .O(N__11087),
            .I(N__11077));
    LocalMux I__1738 (
            .O(N__11084),
            .I(N__11074));
    InMux I__1737 (
            .O(N__11083),
            .I(N__11071));
    InMux I__1736 (
            .O(N__11080),
            .I(N__11068));
    Span4Mux_h I__1735 (
            .O(N__11077),
            .I(N__11063));
    Span4Mux_h I__1734 (
            .O(N__11074),
            .I(N__11063));
    LocalMux I__1733 (
            .O(N__11071),
            .I(N__11058));
    LocalMux I__1732 (
            .O(N__11068),
            .I(N__11058));
    Sp12to4 I__1731 (
            .O(N__11063),
            .I(N__11053));
    Span12Mux_s4_h I__1730 (
            .O(N__11058),
            .I(N__11053));
    Odrv12 I__1729 (
            .O(N__11053),
            .I(\ufifo.txDataValidDZ0 ));
    InMux I__1728 (
            .O(N__11050),
            .I(N__11047));
    LocalMux I__1727 (
            .O(N__11047),
            .I(\ufifo.emitcrlf_fsm.cstate_srsts_sn_1 ));
    CascadeMux I__1726 (
            .O(N__11044),
            .I(\ufifo.N_57_0_1_cascade_ ));
    InMux I__1725 (
            .O(N__11041),
            .I(N__11036));
    InMux I__1724 (
            .O(N__11040),
            .I(N__11033));
    InMux I__1723 (
            .O(N__11039),
            .I(N__11030));
    LocalMux I__1722 (
            .O(N__11036),
            .I(N__11027));
    LocalMux I__1721 (
            .O(N__11033),
            .I(N__11024));
    LocalMux I__1720 (
            .O(N__11030),
            .I(N__11017));
    Span4Mux_h I__1719 (
            .O(N__11027),
            .I(N__11017));
    Span4Mux_h I__1718 (
            .O(N__11024),
            .I(N__11017));
    Odrv4 I__1717 (
            .O(N__11017),
            .I(\Lab_UT.scdp.prng_lfsr_23 ));
    InMux I__1716 (
            .O(N__11014),
            .I(N__11010));
    CascadeMux I__1715 (
            .O(N__11013),
            .I(N__11007));
    LocalMux I__1714 (
            .O(N__11010),
            .I(N__11004));
    InMux I__1713 (
            .O(N__11007),
            .I(N__11001));
    Odrv4 I__1712 (
            .O(N__11004),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24 ));
    LocalMux I__1711 (
            .O(N__11001),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24 ));
    InMux I__1710 (
            .O(N__10996),
            .I(N__10992));
    InMux I__1709 (
            .O(N__10995),
            .I(N__10989));
    LocalMux I__1708 (
            .O(N__10992),
            .I(N__10986));
    LocalMux I__1707 (
            .O(N__10989),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19 ));
    Odrv4 I__1706 (
            .O(N__10986),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19 ));
    InMux I__1705 (
            .O(N__10981),
            .I(N__10977));
    InMux I__1704 (
            .O(N__10980),
            .I(N__10974));
    LocalMux I__1703 (
            .O(N__10977),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20 ));
    LocalMux I__1702 (
            .O(N__10974),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20 ));
    CascadeMux I__1701 (
            .O(N__10969),
            .I(N__10965));
    InMux I__1700 (
            .O(N__10968),
            .I(N__10962));
    InMux I__1699 (
            .O(N__10965),
            .I(N__10959));
    LocalMux I__1698 (
            .O(N__10962),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28 ));
    LocalMux I__1697 (
            .O(N__10959),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28 ));
    InMux I__1696 (
            .O(N__10954),
            .I(N__10951));
    LocalMux I__1695 (
            .O(N__10951),
            .I(N__10946));
    InMux I__1694 (
            .O(N__10950),
            .I(N__10943));
    InMux I__1693 (
            .O(N__10949),
            .I(N__10940));
    Span4Mux_h I__1692 (
            .O(N__10946),
            .I(N__10937));
    LocalMux I__1691 (
            .O(N__10943),
            .I(N__10932));
    LocalMux I__1690 (
            .O(N__10940),
            .I(N__10932));
    Odrv4 I__1689 (
            .O(N__10937),
            .I(\Lab_UT.scdp.prng_lfsr_7 ));
    Odrv4 I__1688 (
            .O(N__10932),
            .I(\Lab_UT.scdp.prng_lfsr_7 ));
    InMux I__1687 (
            .O(N__10927),
            .I(N__10923));
    InMux I__1686 (
            .O(N__10926),
            .I(N__10920));
    LocalMux I__1685 (
            .O(N__10923),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8 ));
    LocalMux I__1684 (
            .O(N__10920),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8 ));
    CascadeMux I__1683 (
            .O(N__10915),
            .I(N__10911));
    InMux I__1682 (
            .O(N__10914),
            .I(N__10908));
    InMux I__1681 (
            .O(N__10911),
            .I(N__10905));
    LocalMux I__1680 (
            .O(N__10908),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26 ));
    LocalMux I__1679 (
            .O(N__10905),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26 ));
    CascadeMux I__1678 (
            .O(N__10900),
            .I(N__10896));
    InMux I__1677 (
            .O(N__10899),
            .I(N__10893));
    InMux I__1676 (
            .O(N__10896),
            .I(N__10890));
    LocalMux I__1675 (
            .O(N__10893),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27 ));
    LocalMux I__1674 (
            .O(N__10890),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27 ));
    InMux I__1673 (
            .O(N__10885),
            .I(N__10881));
    InMux I__1672 (
            .O(N__10884),
            .I(N__10878));
    LocalMux I__1671 (
            .O(N__10881),
            .I(N__10875));
    LocalMux I__1670 (
            .O(N__10878),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21 ));
    Odrv4 I__1669 (
            .O(N__10875),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21 ));
    InMux I__1668 (
            .O(N__10870),
            .I(N__10866));
    CascadeMux I__1667 (
            .O(N__10869),
            .I(N__10863));
    LocalMux I__1666 (
            .O(N__10866),
            .I(N__10860));
    InMux I__1665 (
            .O(N__10863),
            .I(N__10857));
    Odrv4 I__1664 (
            .O(N__10860),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29 ));
    LocalMux I__1663 (
            .O(N__10857),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29 ));
    InMux I__1662 (
            .O(N__10852),
            .I(N__10849));
    LocalMux I__1661 (
            .O(N__10849),
            .I(N__10846));
    Span4Mux_v I__1660 (
            .O(N__10846),
            .I(N__10843));
    Odrv4 I__1659 (
            .O(N__10843),
            .I(\Lab_UT.scdp.d2eData_3_5 ));
    InMux I__1658 (
            .O(N__10840),
            .I(N__10836));
    InMux I__1657 (
            .O(N__10839),
            .I(N__10833));
    LocalMux I__1656 (
            .O(N__10836),
            .I(N__10830));
    LocalMux I__1655 (
            .O(N__10833),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22 ));
    Odrv4 I__1654 (
            .O(N__10830),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22 ));
    InMux I__1653 (
            .O(N__10825),
            .I(N__10821));
    InMux I__1652 (
            .O(N__10824),
            .I(N__10818));
    LocalMux I__1651 (
            .O(N__10821),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18 ));
    LocalMux I__1650 (
            .O(N__10818),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18 ));
    CascadeMux I__1649 (
            .O(N__10813),
            .I(N__10809));
    InMux I__1648 (
            .O(N__10812),
            .I(N__10806));
    InMux I__1647 (
            .O(N__10809),
            .I(N__10803));
    LocalMux I__1646 (
            .O(N__10806),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25 ));
    LocalMux I__1645 (
            .O(N__10803),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25 ));
    InMux I__1644 (
            .O(N__10798),
            .I(N__10794));
    CascadeMux I__1643 (
            .O(N__10797),
            .I(N__10791));
    LocalMux I__1642 (
            .O(N__10794),
            .I(N__10787));
    InMux I__1641 (
            .O(N__10791),
            .I(N__10784));
    InMux I__1640 (
            .O(N__10790),
            .I(N__10781));
    Span4Mux_h I__1639 (
            .O(N__10787),
            .I(N__10778));
    LocalMux I__1638 (
            .O(N__10784),
            .I(N__10775));
    LocalMux I__1637 (
            .O(N__10781),
            .I(\Lab_UT.scdp.prng_lfsr_15 ));
    Odrv4 I__1636 (
            .O(N__10778),
            .I(\Lab_UT.scdp.prng_lfsr_15 ));
    Odrv4 I__1635 (
            .O(N__10775),
            .I(\Lab_UT.scdp.prng_lfsr_15 ));
    InMux I__1634 (
            .O(N__10768),
            .I(N__10764));
    InMux I__1633 (
            .O(N__10767),
            .I(N__10761));
    LocalMux I__1632 (
            .O(N__10764),
            .I(N__10758));
    LocalMux I__1631 (
            .O(N__10761),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16 ));
    Odrv4 I__1630 (
            .O(N__10758),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16 ));
    InMux I__1629 (
            .O(N__10753),
            .I(N__10749));
    InMux I__1628 (
            .O(N__10752),
            .I(N__10746));
    LocalMux I__1627 (
            .O(N__10749),
            .I(N__10743));
    LocalMux I__1626 (
            .O(N__10746),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_3 ));
    Odrv4 I__1625 (
            .O(N__10743),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_3 ));
    InMux I__1624 (
            .O(N__10738),
            .I(N__10734));
    InMux I__1623 (
            .O(N__10737),
            .I(N__10731));
    LocalMux I__1622 (
            .O(N__10734),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9 ));
    LocalMux I__1621 (
            .O(N__10731),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9 ));
    InMux I__1620 (
            .O(N__10726),
            .I(N__10722));
    InMux I__1619 (
            .O(N__10725),
            .I(N__10719));
    LocalMux I__1618 (
            .O(N__10722),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10 ));
    LocalMux I__1617 (
            .O(N__10719),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10 ));
    InMux I__1616 (
            .O(N__10714),
            .I(N__10711));
    LocalMux I__1615 (
            .O(N__10711),
            .I(N__10707));
    InMux I__1614 (
            .O(N__10710),
            .I(N__10704));
    Span4Mux_h I__1613 (
            .O(N__10707),
            .I(N__10701));
    LocalMux I__1612 (
            .O(N__10704),
            .I(N__10698));
    Span4Mux_v I__1611 (
            .O(N__10701),
            .I(N__10695));
    Odrv12 I__1610 (
            .O(N__10698),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    Odrv4 I__1609 (
            .O(N__10695),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    InMux I__1608 (
            .O(N__10690),
            .I(N__10686));
    InMux I__1607 (
            .O(N__10689),
            .I(N__10683));
    LocalMux I__1606 (
            .O(N__10686),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17 ));
    LocalMux I__1605 (
            .O(N__10683),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17 ));
    InMux I__1604 (
            .O(N__10678),
            .I(N__10674));
    InMux I__1603 (
            .O(N__10677),
            .I(N__10671));
    LocalMux I__1602 (
            .O(N__10674),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_14 ));
    LocalMux I__1601 (
            .O(N__10671),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_14 ));
    InMux I__1600 (
            .O(N__10666),
            .I(N__10660));
    InMux I__1599 (
            .O(N__10665),
            .I(N__10660));
    LocalMux I__1598 (
            .O(N__10660),
            .I(\Lab_UT.de_bigL_0 ));
    InMux I__1597 (
            .O(N__10657),
            .I(N__10653));
    InMux I__1596 (
            .O(N__10656),
            .I(N__10644));
    LocalMux I__1595 (
            .O(N__10653),
            .I(N__10641));
    InMux I__1594 (
            .O(N__10652),
            .I(N__10636));
    InMux I__1593 (
            .O(N__10651),
            .I(N__10636));
    InMux I__1592 (
            .O(N__10650),
            .I(N__10633));
    InMux I__1591 (
            .O(N__10649),
            .I(N__10630));
    InMux I__1590 (
            .O(N__10648),
            .I(N__10627));
    InMux I__1589 (
            .O(N__10647),
            .I(N__10624));
    LocalMux I__1588 (
            .O(N__10644),
            .I(buart__rx_bitcount_3));
    Odrv4 I__1587 (
            .O(N__10641),
            .I(buart__rx_bitcount_3));
    LocalMux I__1586 (
            .O(N__10636),
            .I(buart__rx_bitcount_3));
    LocalMux I__1585 (
            .O(N__10633),
            .I(buart__rx_bitcount_3));
    LocalMux I__1584 (
            .O(N__10630),
            .I(buart__rx_bitcount_3));
    LocalMux I__1583 (
            .O(N__10627),
            .I(buart__rx_bitcount_3));
    LocalMux I__1582 (
            .O(N__10624),
            .I(buart__rx_bitcount_3));
    InMux I__1581 (
            .O(N__10609),
            .I(N__10605));
    InMux I__1580 (
            .O(N__10608),
            .I(N__10600));
    LocalMux I__1579 (
            .O(N__10605),
            .I(N__10595));
    InMux I__1578 (
            .O(N__10604),
            .I(N__10592));
    InMux I__1577 (
            .O(N__10603),
            .I(N__10586));
    LocalMux I__1576 (
            .O(N__10600),
            .I(N__10583));
    InMux I__1575 (
            .O(N__10599),
            .I(N__10578));
    InMux I__1574 (
            .O(N__10598),
            .I(N__10578));
    Span4Mux_h I__1573 (
            .O(N__10595),
            .I(N__10573));
    LocalMux I__1572 (
            .O(N__10592),
            .I(N__10573));
    InMux I__1571 (
            .O(N__10591),
            .I(N__10570));
    InMux I__1570 (
            .O(N__10590),
            .I(N__10565));
    InMux I__1569 (
            .O(N__10589),
            .I(N__10565));
    LocalMux I__1568 (
            .O(N__10586),
            .I(buart__rx_bitcount_0));
    Odrv4 I__1567 (
            .O(N__10583),
            .I(buart__rx_bitcount_0));
    LocalMux I__1566 (
            .O(N__10578),
            .I(buart__rx_bitcount_0));
    Odrv4 I__1565 (
            .O(N__10573),
            .I(buart__rx_bitcount_0));
    LocalMux I__1564 (
            .O(N__10570),
            .I(buart__rx_bitcount_0));
    LocalMux I__1563 (
            .O(N__10565),
            .I(buart__rx_bitcount_0));
    InMux I__1562 (
            .O(N__10552),
            .I(N__10541));
    InMux I__1561 (
            .O(N__10551),
            .I(N__10541));
    InMux I__1560 (
            .O(N__10550),
            .I(N__10536));
    InMux I__1559 (
            .O(N__10549),
            .I(N__10536));
    CascadeMux I__1558 (
            .O(N__10548),
            .I(N__10531));
    InMux I__1557 (
            .O(N__10547),
            .I(N__10528));
    InMux I__1556 (
            .O(N__10546),
            .I(N__10525));
    LocalMux I__1555 (
            .O(N__10541),
            .I(N__10522));
    LocalMux I__1554 (
            .O(N__10536),
            .I(N__10519));
    InMux I__1553 (
            .O(N__10535),
            .I(N__10516));
    InMux I__1552 (
            .O(N__10534),
            .I(N__10511));
    InMux I__1551 (
            .O(N__10531),
            .I(N__10511));
    LocalMux I__1550 (
            .O(N__10528),
            .I(buart__rx_bitcount_1));
    LocalMux I__1549 (
            .O(N__10525),
            .I(buart__rx_bitcount_1));
    Odrv4 I__1548 (
            .O(N__10522),
            .I(buart__rx_bitcount_1));
    Odrv4 I__1547 (
            .O(N__10519),
            .I(buart__rx_bitcount_1));
    LocalMux I__1546 (
            .O(N__10516),
            .I(buart__rx_bitcount_1));
    LocalMux I__1545 (
            .O(N__10511),
            .I(buart__rx_bitcount_1));
    CascadeMux I__1544 (
            .O(N__10498),
            .I(N__10491));
    InMux I__1543 (
            .O(N__10497),
            .I(N__10487));
    InMux I__1542 (
            .O(N__10496),
            .I(N__10481));
    InMux I__1541 (
            .O(N__10495),
            .I(N__10481));
    InMux I__1540 (
            .O(N__10494),
            .I(N__10478));
    InMux I__1539 (
            .O(N__10491),
            .I(N__10474));
    InMux I__1538 (
            .O(N__10490),
            .I(N__10471));
    LocalMux I__1537 (
            .O(N__10487),
            .I(N__10468));
    InMux I__1536 (
            .O(N__10486),
            .I(N__10465));
    LocalMux I__1535 (
            .O(N__10481),
            .I(N__10460));
    LocalMux I__1534 (
            .O(N__10478),
            .I(N__10460));
    InMux I__1533 (
            .O(N__10477),
            .I(N__10457));
    LocalMux I__1532 (
            .O(N__10474),
            .I(buart__rx_bitcount_4));
    LocalMux I__1531 (
            .O(N__10471),
            .I(buart__rx_bitcount_4));
    Odrv12 I__1530 (
            .O(N__10468),
            .I(buart__rx_bitcount_4));
    LocalMux I__1529 (
            .O(N__10465),
            .I(buart__rx_bitcount_4));
    Odrv4 I__1528 (
            .O(N__10460),
            .I(buart__rx_bitcount_4));
    LocalMux I__1527 (
            .O(N__10457),
            .I(buart__rx_bitcount_4));
    InMux I__1526 (
            .O(N__10444),
            .I(N__10441));
    LocalMux I__1525 (
            .O(N__10441),
            .I(\buart.Z_rx.shifter_0_fast_RNI1CIH1Z0Z_2 ));
    CascadeMux I__1524 (
            .O(N__10438),
            .I(\buart.Z_rx.bitcount_es_RNIF6D61Z0Z_4_cascade_ ));
    InMux I__1523 (
            .O(N__10435),
            .I(N__10432));
    LocalMux I__1522 (
            .O(N__10432),
            .I(Lab_UT_dk_de_bigD_0));
    InMux I__1521 (
            .O(N__10429),
            .I(N__10426));
    LocalMux I__1520 (
            .O(N__10426),
            .I(\Lab_UT.dk.de_bigD_sxZ0 ));
    CascadeMux I__1519 (
            .O(N__10423),
            .I(Lab_UT_dk_de_bigD_0_cascade_));
    InMux I__1518 (
            .O(N__10420),
            .I(N__10416));
    InMux I__1517 (
            .O(N__10419),
            .I(N__10413));
    LocalMux I__1516 (
            .O(N__10416),
            .I(\Lab_UT.dk.de_bigD_1Z0Z_0 ));
    LocalMux I__1515 (
            .O(N__10413),
            .I(\Lab_UT.dk.de_bigD_1Z0Z_0 ));
    CascadeMux I__1514 (
            .O(N__10408),
            .I(N__10405));
    InMux I__1513 (
            .O(N__10405),
            .I(N__10402));
    LocalMux I__1512 (
            .O(N__10402),
            .I(N__10399));
    Span4Mux_h I__1511 (
            .O(N__10399),
            .I(N__10396));
    Odrv4 I__1510 (
            .O(N__10396),
            .I(\buart.Z_rx.N_41_i_1 ));
    CascadeMux I__1509 (
            .O(N__10393),
            .I(N__10390));
    InMux I__1508 (
            .O(N__10390),
            .I(N__10387));
    LocalMux I__1507 (
            .O(N__10387),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    InMux I__1506 (
            .O(N__10384),
            .I(N__10381));
    LocalMux I__1505 (
            .O(N__10381),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    CascadeMux I__1504 (
            .O(N__10378),
            .I(N__10374));
    InMux I__1503 (
            .O(N__10377),
            .I(N__10368));
    InMux I__1502 (
            .O(N__10374),
            .I(N__10368));
    CascadeMux I__1501 (
            .O(N__10373),
            .I(N__10361));
    LocalMux I__1500 (
            .O(N__10368),
            .I(N__10354));
    InMux I__1499 (
            .O(N__10367),
            .I(N__10351));
    InMux I__1498 (
            .O(N__10366),
            .I(N__10346));
    InMux I__1497 (
            .O(N__10365),
            .I(N__10346));
    InMux I__1496 (
            .O(N__10364),
            .I(N__10343));
    InMux I__1495 (
            .O(N__10361),
            .I(N__10334));
    InMux I__1494 (
            .O(N__10360),
            .I(N__10334));
    InMux I__1493 (
            .O(N__10359),
            .I(N__10334));
    InMux I__1492 (
            .O(N__10358),
            .I(N__10334));
    InMux I__1491 (
            .O(N__10357),
            .I(N__10331));
    Span4Mux_v I__1490 (
            .O(N__10354),
            .I(N__10328));
    LocalMux I__1489 (
            .O(N__10351),
            .I(N__10321));
    LocalMux I__1488 (
            .O(N__10346),
            .I(N__10321));
    LocalMux I__1487 (
            .O(N__10343),
            .I(N__10321));
    LocalMux I__1486 (
            .O(N__10334),
            .I(N__10314));
    LocalMux I__1485 (
            .O(N__10331),
            .I(N__10314));
    Span4Mux_h I__1484 (
            .O(N__10328),
            .I(N__10314));
    Odrv12 I__1483 (
            .O(N__10321),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__1482 (
            .O(N__10314),
            .I(\buart.Z_rx.startbit ));
    InMux I__1481 (
            .O(N__10309),
            .I(N__10296));
    InMux I__1480 (
            .O(N__10308),
            .I(N__10296));
    InMux I__1479 (
            .O(N__10307),
            .I(N__10296));
    InMux I__1478 (
            .O(N__10306),
            .I(N__10296));
    InMux I__1477 (
            .O(N__10305),
            .I(N__10293));
    LocalMux I__1476 (
            .O(N__10296),
            .I(\buart.Z_rx.N_45 ));
    LocalMux I__1475 (
            .O(N__10293),
            .I(\buart.Z_rx.N_45 ));
    CascadeMux I__1474 (
            .O(N__10288),
            .I(N__10285));
    InMux I__1473 (
            .O(N__10285),
            .I(N__10282));
    LocalMux I__1472 (
            .O(N__10282),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    CEMux I__1471 (
            .O(N__10279),
            .I(N__10275));
    CEMux I__1470 (
            .O(N__10278),
            .I(N__10272));
    LocalMux I__1469 (
            .O(N__10275),
            .I(N__10269));
    LocalMux I__1468 (
            .O(N__10272),
            .I(N__10266));
    Span4Mux_v I__1467 (
            .O(N__10269),
            .I(N__10263));
    Odrv4 I__1466 (
            .O(N__10266),
            .I(\buart.Z_rx.N_43 ));
    Odrv4 I__1465 (
            .O(N__10263),
            .I(\buart.Z_rx.N_43 ));
    CascadeMux I__1464 (
            .O(N__10258),
            .I(N__10255));
    InMux I__1463 (
            .O(N__10255),
            .I(N__10252));
    LocalMux I__1462 (
            .O(N__10252),
            .I(\Lab_UT.dk.de_bigL_sxZ0 ));
    InMux I__1461 (
            .O(N__10249),
            .I(N__10246));
    LocalMux I__1460 (
            .O(N__10246),
            .I(\Lab_UT.de_bigL_3 ));
    InMux I__1459 (
            .O(N__10243),
            .I(N__10240));
    LocalMux I__1458 (
            .O(N__10240),
            .I(N__10237));
    Odrv4 I__1457 (
            .O(N__10237),
            .I(\Lab_UT.scctrl.g0_17_N_3LZ0Z3 ));
    CascadeMux I__1456 (
            .O(N__10234),
            .I(\Lab_UT.de_bigL_3_cascade_ ));
    InMux I__1455 (
            .O(N__10231),
            .I(N__10228));
    LocalMux I__1454 (
            .O(N__10228),
            .I(N__10225));
    Odrv4 I__1453 (
            .O(N__10225),
            .I(\Lab_UT.scctrl.g0_17_N_2LZ0Z1 ));
    CascadeMux I__1452 (
            .O(N__10222),
            .I(\buart.Z_rx.N_58_cascade_ ));
    InMux I__1451 (
            .O(N__10219),
            .I(N__10216));
    LocalMux I__1450 (
            .O(N__10216),
            .I(N__10213));
    Span4Mux_h I__1449 (
            .O(N__10213),
            .I(N__10209));
    InMux I__1448 (
            .O(N__10212),
            .I(N__10206));
    Span4Mux_v I__1447 (
            .O(N__10209),
            .I(N__10203));
    LocalMux I__1446 (
            .O(N__10206),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    Odrv4 I__1445 (
            .O(N__10203),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    InMux I__1444 (
            .O(N__10198),
            .I(N__10194));
    InMux I__1443 (
            .O(N__10197),
            .I(N__10191));
    LocalMux I__1442 (
            .O(N__10194),
            .I(\buart.Z_rx.N_58 ));
    LocalMux I__1441 (
            .O(N__10191),
            .I(\buart.Z_rx.N_58 ));
    CascadeMux I__1440 (
            .O(N__10186),
            .I(\buart.Z_rx.startbit_cascade_ ));
    InMux I__1439 (
            .O(N__10183),
            .I(N__10179));
    CascadeMux I__1438 (
            .O(N__10182),
            .I(N__10175));
    LocalMux I__1437 (
            .O(N__10179),
            .I(N__10172));
    InMux I__1436 (
            .O(N__10178),
            .I(N__10167));
    InMux I__1435 (
            .O(N__10175),
            .I(N__10164));
    Span4Mux_h I__1434 (
            .O(N__10172),
            .I(N__10161));
    InMux I__1433 (
            .O(N__10171),
            .I(N__10156));
    InMux I__1432 (
            .O(N__10170),
            .I(N__10156));
    LocalMux I__1431 (
            .O(N__10167),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__1430 (
            .O(N__10164),
            .I(\buart.Z_rx.ser_clk ));
    Odrv4 I__1429 (
            .O(N__10161),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__1428 (
            .O(N__10156),
            .I(\buart.Z_rx.ser_clk ));
    InMux I__1427 (
            .O(N__10147),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__1426 (
            .O(N__10144),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    InMux I__1425 (
            .O(N__10141),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__1424 (
            .O(N__10138),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    CascadeMux I__1423 (
            .O(N__10135),
            .I(N__10131));
    InMux I__1422 (
            .O(N__10134),
            .I(N__10128));
    InMux I__1421 (
            .O(N__10131),
            .I(N__10125));
    LocalMux I__1420 (
            .O(N__10128),
            .I(N__10122));
    LocalMux I__1419 (
            .O(N__10125),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    Odrv4 I__1418 (
            .O(N__10122),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__1417 (
            .O(N__10117),
            .I(N__10113));
    InMux I__1416 (
            .O(N__10116),
            .I(N__10110));
    InMux I__1415 (
            .O(N__10113),
            .I(N__10107));
    LocalMux I__1414 (
            .O(N__10110),
            .I(N__10104));
    LocalMux I__1413 (
            .O(N__10107),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    Odrv4 I__1412 (
            .O(N__10104),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    CascadeMux I__1411 (
            .O(N__10099),
            .I(N__10096));
    InMux I__1410 (
            .O(N__10096),
            .I(N__10092));
    InMux I__1409 (
            .O(N__10095),
            .I(N__10089));
    LocalMux I__1408 (
            .O(N__10092),
            .I(N__10086));
    LocalMux I__1407 (
            .O(N__10089),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    Odrv12 I__1406 (
            .O(N__10086),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    InMux I__1405 (
            .O(N__10081),
            .I(N__10078));
    LocalMux I__1404 (
            .O(N__10078),
            .I(\ufifo.fifo.un1_emptyB_NE_2 ));
    InMux I__1403 (
            .O(N__10075),
            .I(N__10072));
    LocalMux I__1402 (
            .O(N__10072),
            .I(N__10069));
    Odrv4 I__1401 (
            .O(N__10069),
            .I(\ufifo.fifo.un1_emptyB_NE_1 ));
    CascadeMux I__1400 (
            .O(N__10066),
            .I(N__10063));
    InMux I__1399 (
            .O(N__10063),
            .I(N__10060));
    LocalMux I__1398 (
            .O(N__10060),
            .I(N__10057));
    Odrv4 I__1397 (
            .O(N__10057),
            .I(\ufifo.fifo.un1_emptyB_NE_3 ));
    InMux I__1396 (
            .O(N__10054),
            .I(N__10051));
    LocalMux I__1395 (
            .O(N__10051),
            .I(N__10048));
    Odrv4 I__1394 (
            .O(N__10048),
            .I(\ufifo.fifo.un1_emptyB_NE_4 ));
    CascadeMux I__1393 (
            .O(N__10045),
            .I(\ufifo.emptyB_0_cascade_ ));
    CascadeMux I__1392 (
            .O(N__10042),
            .I(N__10039));
    InMux I__1391 (
            .O(N__10039),
            .I(N__10033));
    InMux I__1390 (
            .O(N__10038),
            .I(N__10033));
    LocalMux I__1389 (
            .O(N__10033),
            .I(\ufifo.tx_fsm.cstateZ0Z_1 ));
    CascadeMux I__1388 (
            .O(N__10030),
            .I(\ufifo.tx_fsm.N_62_0_cascade_ ));
    CascadeMux I__1387 (
            .O(N__10027),
            .I(N__10020));
    SRMux I__1386 (
            .O(N__10026),
            .I(N__10017));
    CEMux I__1385 (
            .O(N__10025),
            .I(N__10014));
    InMux I__1384 (
            .O(N__10024),
            .I(N__10011));
    InMux I__1383 (
            .O(N__10023),
            .I(N__10008));
    InMux I__1382 (
            .O(N__10020),
            .I(N__10005));
    LocalMux I__1381 (
            .O(N__10017),
            .I(N__10002));
    LocalMux I__1380 (
            .O(N__10014),
            .I(N__9999));
    LocalMux I__1379 (
            .O(N__10011),
            .I(N__9996));
    LocalMux I__1378 (
            .O(N__10008),
            .I(N__9991));
    LocalMux I__1377 (
            .O(N__10005),
            .I(N__9991));
    Span4Mux_h I__1376 (
            .O(N__10002),
            .I(N__9988));
    Span4Mux_h I__1375 (
            .O(N__9999),
            .I(N__9985));
    Span4Mux_h I__1374 (
            .O(N__9996),
            .I(N__9980));
    Span4Mux_s2_v I__1373 (
            .O(N__9991),
            .I(N__9980));
    Odrv4 I__1372 (
            .O(N__9988),
            .I(\ufifo.popFifo ));
    Odrv4 I__1371 (
            .O(N__9985),
            .I(\ufifo.popFifo ));
    Odrv4 I__1370 (
            .O(N__9980),
            .I(\ufifo.popFifo ));
    SRMux I__1369 (
            .O(N__9973),
            .I(N__9970));
    LocalMux I__1368 (
            .O(N__9970),
            .I(N__9967));
    Span4Mux_v I__1367 (
            .O(N__9967),
            .I(N__9963));
    SRMux I__1366 (
            .O(N__9966),
            .I(N__9960));
    Sp12to4 I__1365 (
            .O(N__9963),
            .I(N__9956));
    LocalMux I__1364 (
            .O(N__9960),
            .I(N__9953));
    SRMux I__1363 (
            .O(N__9959),
            .I(N__9950));
    Odrv12 I__1362 (
            .O(N__9956),
            .I(rst_i_3_i));
    Odrv4 I__1361 (
            .O(N__9953),
            .I(rst_i_3_i));
    LocalMux I__1360 (
            .O(N__9950),
            .I(rst_i_3_i));
    InMux I__1359 (
            .O(N__9943),
            .I(N__9938));
    InMux I__1358 (
            .O(N__9942),
            .I(N__9935));
    InMux I__1357 (
            .O(N__9941),
            .I(N__9932));
    LocalMux I__1356 (
            .O(N__9938),
            .I(N__9928));
    LocalMux I__1355 (
            .O(N__9935),
            .I(N__9925));
    LocalMux I__1354 (
            .O(N__9932),
            .I(N__9921));
    CascadeMux I__1353 (
            .O(N__9931),
            .I(N__9918));
    Span4Mux_v I__1352 (
            .O(N__9928),
            .I(N__9911));
    Span4Mux_v I__1351 (
            .O(N__9925),
            .I(N__9911));
    InMux I__1350 (
            .O(N__9924),
            .I(N__9908));
    Span4Mux_v I__1349 (
            .O(N__9921),
            .I(N__9905));
    InMux I__1348 (
            .O(N__9918),
            .I(N__9900));
    InMux I__1347 (
            .O(N__9917),
            .I(N__9900));
    InMux I__1346 (
            .O(N__9916),
            .I(N__9897));
    Span4Mux_h I__1345 (
            .O(N__9911),
            .I(N__9892));
    LocalMux I__1344 (
            .O(N__9908),
            .I(N__9892));
    Odrv4 I__1343 (
            .O(N__9905),
            .I(\ufifo.emitcrlf_fsm.cstateZ0Z_0 ));
    LocalMux I__1342 (
            .O(N__9900),
            .I(\ufifo.emitcrlf_fsm.cstateZ0Z_0 ));
    LocalMux I__1341 (
            .O(N__9897),
            .I(\ufifo.emitcrlf_fsm.cstateZ0Z_0 ));
    Odrv4 I__1340 (
            .O(N__9892),
            .I(\ufifo.emitcrlf_fsm.cstateZ0Z_0 ));
    CascadeMux I__1339 (
            .O(N__9883),
            .I(\buart.Z_rx.bitcountlde_i_o2_0_cascade_ ));
    InMux I__1338 (
            .O(N__9880),
            .I(N__9877));
    LocalMux I__1337 (
            .O(N__9877),
            .I(N__9874));
    Odrv12 I__1336 (
            .O(N__9874),
            .I(\Lab_UT.scdp.lsBitsi.q_esr_RNI0TMAZ0Z_3 ));
    CascadeMux I__1335 (
            .O(N__9871),
            .I(\Lab_UT.scdp.q_RNIRM8BD_3_cascade_ ));
    InMux I__1334 (
            .O(N__9868),
            .I(N__9865));
    LocalMux I__1333 (
            .O(N__9865),
            .I(N__9862));
    Span4Mux_s3_h I__1332 (
            .O(N__9862),
            .I(N__9859));
    Span4Mux_v I__1331 (
            .O(N__9859),
            .I(N__9856));
    Odrv4 I__1330 (
            .O(N__9856),
            .I(\ufifo.txdataDZ0Z_3 ));
    InMux I__1329 (
            .O(N__9853),
            .I(N__9850));
    LocalMux I__1328 (
            .O(N__9850),
            .I(N__9845));
    InMux I__1327 (
            .O(N__9849),
            .I(N__9842));
    InMux I__1326 (
            .O(N__9848),
            .I(N__9839));
    Span12Mux_s10_v I__1325 (
            .O(N__9845),
            .I(N__9836));
    LocalMux I__1324 (
            .O(N__9842),
            .I(N__9833));
    LocalMux I__1323 (
            .O(N__9839),
            .I(\Lab_UT.scdp.byteToDecrypt_0 ));
    Odrv12 I__1322 (
            .O(N__9836),
            .I(\Lab_UT.scdp.byteToDecrypt_0 ));
    Odrv4 I__1321 (
            .O(N__9833),
            .I(\Lab_UT.scdp.byteToDecrypt_0 ));
    InMux I__1320 (
            .O(N__9826),
            .I(N__9821));
    InMux I__1319 (
            .O(N__9825),
            .I(N__9818));
    InMux I__1318 (
            .O(N__9824),
            .I(N__9815));
    LocalMux I__1317 (
            .O(N__9821),
            .I(\Lab_UT.scdp.byteToDecrypt_3 ));
    LocalMux I__1316 (
            .O(N__9818),
            .I(\Lab_UT.scdp.byteToDecrypt_3 ));
    LocalMux I__1315 (
            .O(N__9815),
            .I(\Lab_UT.scdp.byteToDecrypt_3 ));
    CascadeMux I__1314 (
            .O(N__9808),
            .I(N__9805));
    InMux I__1313 (
            .O(N__9805),
            .I(N__9802));
    LocalMux I__1312 (
            .O(N__9802),
            .I(N__9799));
    Span4Mux_v I__1311 (
            .O(N__9799),
            .I(N__9794));
    InMux I__1310 (
            .O(N__9798),
            .I(N__9791));
    InMux I__1309 (
            .O(N__9797),
            .I(N__9788));
    Odrv4 I__1308 (
            .O(N__9794),
            .I(\ufifo.fifo.wraddrZ0Z_4 ));
    LocalMux I__1307 (
            .O(N__9791),
            .I(\ufifo.fifo.wraddrZ0Z_4 ));
    LocalMux I__1306 (
            .O(N__9788),
            .I(\ufifo.fifo.wraddrZ0Z_4 ));
    CascadeMux I__1305 (
            .O(N__9781),
            .I(N__9778));
    InMux I__1304 (
            .O(N__9778),
            .I(N__9775));
    LocalMux I__1303 (
            .O(N__9775),
            .I(N__9771));
    InMux I__1302 (
            .O(N__9774),
            .I(N__9767));
    Span4Mux_v I__1301 (
            .O(N__9771),
            .I(N__9764));
    InMux I__1300 (
            .O(N__9770),
            .I(N__9761));
    LocalMux I__1299 (
            .O(N__9767),
            .I(N__9758));
    Odrv4 I__1298 (
            .O(N__9764),
            .I(\ufifo.fifo.rdaddrZ0Z_4 ));
    LocalMux I__1297 (
            .O(N__9761),
            .I(\ufifo.fifo.rdaddrZ0Z_4 ));
    Odrv4 I__1296 (
            .O(N__9758),
            .I(\ufifo.fifo.rdaddrZ0Z_4 ));
    CascadeMux I__1295 (
            .O(N__9751),
            .I(N__9748));
    InMux I__1294 (
            .O(N__9748),
            .I(N__9745));
    LocalMux I__1293 (
            .O(N__9745),
            .I(N__9741));
    CascadeMux I__1292 (
            .O(N__9744),
            .I(N__9737));
    Span4Mux_v I__1291 (
            .O(N__9741),
            .I(N__9734));
    InMux I__1290 (
            .O(N__9740),
            .I(N__9731));
    InMux I__1289 (
            .O(N__9737),
            .I(N__9728));
    Odrv4 I__1288 (
            .O(N__9734),
            .I(\ufifo.fifo.wraddrZ0Z_5 ));
    LocalMux I__1287 (
            .O(N__9731),
            .I(\ufifo.fifo.wraddrZ0Z_5 ));
    LocalMux I__1286 (
            .O(N__9728),
            .I(\ufifo.fifo.wraddrZ0Z_5 ));
    CascadeMux I__1285 (
            .O(N__9721),
            .I(N__9718));
    InMux I__1284 (
            .O(N__9718),
            .I(N__9715));
    LocalMux I__1283 (
            .O(N__9715),
            .I(N__9711));
    InMux I__1282 (
            .O(N__9714),
            .I(N__9707));
    Span12Mux_v I__1281 (
            .O(N__9711),
            .I(N__9704));
    InMux I__1280 (
            .O(N__9710),
            .I(N__9701));
    LocalMux I__1279 (
            .O(N__9707),
            .I(N__9698));
    Odrv12 I__1278 (
            .O(N__9704),
            .I(\ufifo.fifo.rdaddrZ0Z_5 ));
    LocalMux I__1277 (
            .O(N__9701),
            .I(\ufifo.fifo.rdaddrZ0Z_5 ));
    Odrv4 I__1276 (
            .O(N__9698),
            .I(\ufifo.fifo.rdaddrZ0Z_5 ));
    CascadeMux I__1275 (
            .O(N__9691),
            .I(N__9688));
    InMux I__1274 (
            .O(N__9688),
            .I(N__9685));
    LocalMux I__1273 (
            .O(N__9685),
            .I(N__9682));
    Span4Mux_v I__1272 (
            .O(N__9682),
            .I(N__9677));
    InMux I__1271 (
            .O(N__9681),
            .I(N__9674));
    InMux I__1270 (
            .O(N__9680),
            .I(N__9671));
    Odrv4 I__1269 (
            .O(N__9677),
            .I(\ufifo.fifo.wraddrZ0Z_2 ));
    LocalMux I__1268 (
            .O(N__9674),
            .I(\ufifo.fifo.wraddrZ0Z_2 ));
    LocalMux I__1267 (
            .O(N__9671),
            .I(\ufifo.fifo.wraddrZ0Z_2 ));
    CascadeMux I__1266 (
            .O(N__9664),
            .I(N__9661));
    InMux I__1265 (
            .O(N__9661),
            .I(N__9658));
    LocalMux I__1264 (
            .O(N__9658),
            .I(N__9654));
    InMux I__1263 (
            .O(N__9657),
            .I(N__9650));
    Span4Mux_v I__1262 (
            .O(N__9654),
            .I(N__9647));
    InMux I__1261 (
            .O(N__9653),
            .I(N__9644));
    LocalMux I__1260 (
            .O(N__9650),
            .I(N__9641));
    Odrv4 I__1259 (
            .O(N__9647),
            .I(\ufifo.fifo.rdaddrZ0Z_3 ));
    LocalMux I__1258 (
            .O(N__9644),
            .I(\ufifo.fifo.rdaddrZ0Z_3 ));
    Odrv4 I__1257 (
            .O(N__9641),
            .I(\ufifo.fifo.rdaddrZ0Z_3 ));
    CascadeMux I__1256 (
            .O(N__9634),
            .I(N__9631));
    InMux I__1255 (
            .O(N__9631),
            .I(N__9628));
    LocalMux I__1254 (
            .O(N__9628),
            .I(N__9624));
    CascadeMux I__1253 (
            .O(N__9627),
            .I(N__9620));
    Span4Mux_v I__1252 (
            .O(N__9624),
            .I(N__9617));
    InMux I__1251 (
            .O(N__9623),
            .I(N__9614));
    InMux I__1250 (
            .O(N__9620),
            .I(N__9611));
    Odrv4 I__1249 (
            .O(N__9617),
            .I(\ufifo.fifo.wraddrZ0Z_3 ));
    LocalMux I__1248 (
            .O(N__9614),
            .I(\ufifo.fifo.wraddrZ0Z_3 ));
    LocalMux I__1247 (
            .O(N__9611),
            .I(\ufifo.fifo.wraddrZ0Z_3 ));
    CascadeMux I__1246 (
            .O(N__9604),
            .I(N__9601));
    InMux I__1245 (
            .O(N__9601),
            .I(N__9598));
    LocalMux I__1244 (
            .O(N__9598),
            .I(N__9594));
    InMux I__1243 (
            .O(N__9597),
            .I(N__9590));
    Span4Mux_v I__1242 (
            .O(N__9594),
            .I(N__9587));
    InMux I__1241 (
            .O(N__9593),
            .I(N__9584));
    LocalMux I__1240 (
            .O(N__9590),
            .I(N__9581));
    Odrv4 I__1239 (
            .O(N__9587),
            .I(\ufifo.fifo.rdaddrZ0Z_2 ));
    LocalMux I__1238 (
            .O(N__9584),
            .I(\ufifo.fifo.rdaddrZ0Z_2 ));
    Odrv4 I__1237 (
            .O(N__9581),
            .I(\ufifo.fifo.rdaddrZ0Z_2 ));
    CascadeMux I__1236 (
            .O(N__9574),
            .I(N__9571));
    InMux I__1235 (
            .O(N__9571),
            .I(N__9568));
    LocalMux I__1234 (
            .O(N__9568),
            .I(N__9563));
    InMux I__1233 (
            .O(N__9567),
            .I(N__9560));
    InMux I__1232 (
            .O(N__9566),
            .I(N__9557));
    Span4Mux_v I__1231 (
            .O(N__9563),
            .I(N__9550));
    LocalMux I__1230 (
            .O(N__9560),
            .I(N__9550));
    LocalMux I__1229 (
            .O(N__9557),
            .I(N__9550));
    Odrv4 I__1228 (
            .O(N__9550),
            .I(\ufifo.fifo.wraddrZ0Z_1 ));
    CascadeMux I__1227 (
            .O(N__9547),
            .I(\ufifo.fifo.un1_emptyB_NE_0_cascade_ ));
    CascadeMux I__1226 (
            .O(N__9544),
            .I(N__9541));
    InMux I__1225 (
            .O(N__9541),
            .I(N__9538));
    LocalMux I__1224 (
            .O(N__9538),
            .I(N__9534));
    InMux I__1223 (
            .O(N__9537),
            .I(N__9531));
    Span4Mux_v I__1222 (
            .O(N__9534),
            .I(N__9527));
    LocalMux I__1221 (
            .O(N__9531),
            .I(N__9524));
    InMux I__1220 (
            .O(N__9530),
            .I(N__9521));
    Span4Mux_v I__1219 (
            .O(N__9527),
            .I(N__9516));
    Span4Mux_h I__1218 (
            .O(N__9524),
            .I(N__9516));
    LocalMux I__1217 (
            .O(N__9521),
            .I(\ufifo.fifo.rdaddrZ0Z_1 ));
    Odrv4 I__1216 (
            .O(N__9516),
            .I(\ufifo.fifo.rdaddrZ0Z_1 ));
    InMux I__1215 (
            .O(N__9511),
            .I(N__9507));
    CascadeMux I__1214 (
            .O(N__9510),
            .I(N__9504));
    LocalMux I__1213 (
            .O(N__9507),
            .I(N__9501));
    InMux I__1212 (
            .O(N__9504),
            .I(N__9498));
    Span4Mux_h I__1211 (
            .O(N__9501),
            .I(N__9495));
    LocalMux I__1210 (
            .O(N__9498),
            .I(N__9492));
    Odrv4 I__1209 (
            .O(N__9495),
            .I(\ufifo.tx_fsm.fifo_txdata_rdy ));
    Odrv12 I__1208 (
            .O(N__9492),
            .I(\ufifo.tx_fsm.fifo_txdata_rdy ));
    InMux I__1207 (
            .O(N__9487),
            .I(N__9484));
    LocalMux I__1206 (
            .O(N__9484),
            .I(N__9480));
    InMux I__1205 (
            .O(N__9483),
            .I(N__9477));
    Odrv4 I__1204 (
            .O(N__9480),
            .I(\Lab_UT.scdp.e2dData_2 ));
    LocalMux I__1203 (
            .O(N__9477),
            .I(\Lab_UT.scdp.e2dData_2 ));
    InMux I__1202 (
            .O(N__9472),
            .I(N__9468));
    InMux I__1201 (
            .O(N__9471),
            .I(N__9465));
    LocalMux I__1200 (
            .O(N__9468),
            .I(\Lab_UT.scdp.N_59_i ));
    LocalMux I__1199 (
            .O(N__9465),
            .I(\Lab_UT.scdp.N_59_i ));
    InMux I__1198 (
            .O(N__9460),
            .I(N__9457));
    LocalMux I__1197 (
            .O(N__9457),
            .I(\Lab_UT.scdp.pinst0.un12_pValidZ0Z_1 ));
    InMux I__1196 (
            .O(N__9454),
            .I(N__9451));
    LocalMux I__1195 (
            .O(N__9451),
            .I(N__9448));
    Odrv12 I__1194 (
            .O(N__9448),
            .I(\Lab_UT.scdp.msBitsi.msBitsD_4 ));
    InMux I__1193 (
            .O(N__9445),
            .I(N__9439));
    InMux I__1192 (
            .O(N__9444),
            .I(N__9439));
    LocalMux I__1191 (
            .O(N__9439),
            .I(N__9435));
    InMux I__1190 (
            .O(N__9438),
            .I(N__9432));
    Odrv12 I__1189 (
            .O(N__9435),
            .I(\Lab_UT.scdp.d2eData_3_4 ));
    LocalMux I__1188 (
            .O(N__9432),
            .I(\Lab_UT.scdp.d2eData_3_4 ));
    CascadeMux I__1187 (
            .O(N__9427),
            .I(\Lab_UT.scdp.d2eData_3_4_cascade_ ));
    CascadeMux I__1186 (
            .O(N__9424),
            .I(\Lab_UT.scdp.q_RNIIAV0D_0_cascade_ ));
    InMux I__1185 (
            .O(N__9421),
            .I(N__9418));
    LocalMux I__1184 (
            .O(N__9418),
            .I(\Lab_UT.scdp.msBitsi.q_esr_RNI239EZ0Z_4 ));
    InMux I__1183 (
            .O(N__9415),
            .I(N__9412));
    LocalMux I__1182 (
            .O(N__9412),
            .I(N__9409));
    Span4Mux_v I__1181 (
            .O(N__9409),
            .I(N__9406));
    Odrv4 I__1180 (
            .O(N__9406),
            .I(\ufifo.txdataDZ0Z_4 ));
    InMux I__1179 (
            .O(N__9403),
            .I(N__9394));
    InMux I__1178 (
            .O(N__9402),
            .I(N__9394));
    InMux I__1177 (
            .O(N__9401),
            .I(N__9394));
    LocalMux I__1176 (
            .O(N__9394),
            .I(N__9390));
    InMux I__1175 (
            .O(N__9393),
            .I(N__9387));
    Odrv4 I__1174 (
            .O(N__9390),
            .I(\Lab_UT.scdp.d2eData_3_3 ));
    LocalMux I__1173 (
            .O(N__9387),
            .I(\Lab_UT.scdp.d2eData_3_3 ));
    InMux I__1172 (
            .O(N__9382),
            .I(N__9376));
    InMux I__1171 (
            .O(N__9381),
            .I(N__9367));
    InMux I__1170 (
            .O(N__9380),
            .I(N__9367));
    InMux I__1169 (
            .O(N__9379),
            .I(N__9367));
    LocalMux I__1168 (
            .O(N__9376),
            .I(N__9364));
    InMux I__1167 (
            .O(N__9375),
            .I(N__9359));
    InMux I__1166 (
            .O(N__9374),
            .I(N__9359));
    LocalMux I__1165 (
            .O(N__9367),
            .I(N__9356));
    Odrv12 I__1164 (
            .O(N__9364),
            .I(\Lab_UT.scdp.pValid_0 ));
    LocalMux I__1163 (
            .O(N__9359),
            .I(\Lab_UT.scdp.pValid_0 ));
    Odrv4 I__1162 (
            .O(N__9356),
            .I(\Lab_UT.scdp.pValid_0 ));
    CascadeMux I__1161 (
            .O(N__9349),
            .I(\Lab_UT.scdp.d2eData_3_3_cascade_ ));
    CascadeMux I__1160 (
            .O(N__9346),
            .I(\Lab_UT.scdp.d2eData_3_2_cascade_ ));
    InMux I__1159 (
            .O(N__9343),
            .I(N__9340));
    LocalMux I__1158 (
            .O(N__9340),
            .I(N__9337));
    Span4Mux_h I__1157 (
            .O(N__9337),
            .I(N__9334));
    Odrv4 I__1156 (
            .O(N__9334),
            .I(\Lab_UT.scdp.u2.byteToEncrypt_2 ));
    CascadeMux I__1155 (
            .O(N__9331),
            .I(N__9328));
    InMux I__1154 (
            .O(N__9328),
            .I(N__9319));
    InMux I__1153 (
            .O(N__9327),
            .I(N__9319));
    InMux I__1152 (
            .O(N__9326),
            .I(N__9319));
    LocalMux I__1151 (
            .O(N__9319),
            .I(\Lab_UT.scdp.d2eData_2 ));
    CascadeMux I__1150 (
            .O(N__9316),
            .I(N__9312));
    InMux I__1149 (
            .O(N__9315),
            .I(N__9304));
    InMux I__1148 (
            .O(N__9312),
            .I(N__9304));
    InMux I__1147 (
            .O(N__9311),
            .I(N__9304));
    LocalMux I__1146 (
            .O(N__9304),
            .I(\Lab_UT.scdp.d2eData_1 ));
    CascadeMux I__1145 (
            .O(N__9301),
            .I(N__9298));
    InMux I__1144 (
            .O(N__9298),
            .I(N__9295));
    LocalMux I__1143 (
            .O(N__9295),
            .I(\Lab_UT.scdp.lsBitsD_2 ));
    InMux I__1142 (
            .O(N__9292),
            .I(N__9288));
    InMux I__1141 (
            .O(N__9291),
            .I(N__9285));
    LocalMux I__1140 (
            .O(N__9288),
            .I(N__9282));
    LocalMux I__1139 (
            .O(N__9285),
            .I(\Lab_UT.scdp.d2eData_3_1 ));
    Odrv4 I__1138 (
            .O(N__9282),
            .I(\Lab_UT.scdp.d2eData_3_1 ));
    CascadeMux I__1137 (
            .O(N__9277),
            .I(\Lab_UT.scdp.pinst0.un12_pValidZ0Z_0_cascade_ ));
    CascadeMux I__1136 (
            .O(N__9274),
            .I(\Lab_UT.scdp.un12_pValid_cascade_ ));
    InMux I__1135 (
            .O(N__9271),
            .I(N__9267));
    InMux I__1134 (
            .O(N__9270),
            .I(N__9264));
    LocalMux I__1133 (
            .O(N__9267),
            .I(N__9261));
    LocalMux I__1132 (
            .O(N__9264),
            .I(N__9258));
    Span12Mux_s11_v I__1131 (
            .O(N__9261),
            .I(N__9254));
    Span4Mux_s3_h I__1130 (
            .O(N__9258),
            .I(N__9251));
    InMux I__1129 (
            .O(N__9257),
            .I(N__9248));
    Odrv12 I__1128 (
            .O(N__9254),
            .I(\Lab_UT.scdp.d2eData_3_0 ));
    Odrv4 I__1127 (
            .O(N__9251),
            .I(\Lab_UT.scdp.d2eData_3_0 ));
    LocalMux I__1126 (
            .O(N__9248),
            .I(\Lab_UT.scdp.d2eData_3_0 ));
    InMux I__1125 (
            .O(N__9241),
            .I(N__9238));
    LocalMux I__1124 (
            .O(N__9238),
            .I(\Lab_UT.scdp.un12_pValid ));
    InMux I__1123 (
            .O(N__9235),
            .I(N__9229));
    InMux I__1122 (
            .O(N__9234),
            .I(N__9229));
    LocalMux I__1121 (
            .O(N__9229),
            .I(N__9226));
    Odrv12 I__1120 (
            .O(N__9226),
            .I(\Lab_UT.scdp.e2dData_6 ));
    InMux I__1119 (
            .O(N__9223),
            .I(N__9220));
    LocalMux I__1118 (
            .O(N__9220),
            .I(N__9217));
    Odrv12 I__1117 (
            .O(N__9217),
            .I(\Lab_UT.scdp.q_RNIDHFGA_3 ));
    InMux I__1116 (
            .O(N__9214),
            .I(N__9211));
    LocalMux I__1115 (
            .O(N__9211),
            .I(\Lab_UT.scdp.d2eData_3_2 ));
    InMux I__1114 (
            .O(N__9208),
            .I(N__9205));
    LocalMux I__1113 (
            .O(N__9205),
            .I(N__9202));
    Span4Mux_v I__1112 (
            .O(N__9202),
            .I(N__9199));
    Odrv4 I__1111 (
            .O(N__9199),
            .I(\Lab_UT.scdp.msBitsi.msBitsD_2 ));
    CascadeMux I__1110 (
            .O(N__9196),
            .I(\Lab_UT.scdp.msBitsi.L4_tx_data_ns_1_2_cascade_ ));
    InMux I__1109 (
            .O(N__9193),
            .I(N__9190));
    LocalMux I__1108 (
            .O(N__9190),
            .I(N__9187));
    Span4Mux_s3_h I__1107 (
            .O(N__9187),
            .I(N__9184));
    Odrv4 I__1106 (
            .O(N__9184),
            .I(\ufifo.txdataDZ0Z_2 ));
    CascadeMux I__1105 (
            .O(N__9181),
            .I(\Lab_UT.scdp.d2eData_3_1_cascade_ ));
    InMux I__1104 (
            .O(N__9178),
            .I(N__9175));
    LocalMux I__1103 (
            .O(N__9175),
            .I(\Lab_UT.scdp.q_RNIABC1D_1 ));
    InMux I__1102 (
            .O(N__9172),
            .I(N__9169));
    LocalMux I__1101 (
            .O(N__9169),
            .I(N__9166));
    Span4Mux_h I__1100 (
            .O(N__9166),
            .I(N__9163));
    Odrv4 I__1099 (
            .O(N__9163),
            .I(\Lab_UT.scdp.u2.byteToEncrypt_1 ));
    CascadeMux I__1098 (
            .O(N__9160),
            .I(\Lab_UT.scdp.d2eData_1_cascade_ ));
    CascadeMux I__1097 (
            .O(N__9157),
            .I(\Lab_UT.scdp.lsBits_6_cascade_ ));
    InMux I__1096 (
            .O(N__9154),
            .I(N__9151));
    LocalMux I__1095 (
            .O(N__9151),
            .I(\Lab_UT.scdp.lsBitsD_1 ));
    InMux I__1094 (
            .O(N__9148),
            .I(N__9145));
    LocalMux I__1093 (
            .O(N__9145),
            .I(N__9142));
    Odrv12 I__1092 (
            .O(N__9142),
            .I(\Lab_UT.scdp.lsBitsi.lsBitsD_3 ));
    InMux I__1091 (
            .O(N__9139),
            .I(N__9130));
    InMux I__1090 (
            .O(N__9138),
            .I(N__9130));
    InMux I__1089 (
            .O(N__9137),
            .I(N__9130));
    LocalMux I__1088 (
            .O(N__9130),
            .I(N__9127));
    Span4Mux_h I__1087 (
            .O(N__9127),
            .I(N__9124));
    Odrv4 I__1086 (
            .O(N__9124),
            .I(\Lab_UT.scdp.byteToEncrypt_3 ));
    InMux I__1085 (
            .O(N__9121),
            .I(N__9118));
    LocalMux I__1084 (
            .O(N__9118),
            .I(N__9115));
    Span4Mux_v I__1083 (
            .O(N__9115),
            .I(N__9112));
    Odrv4 I__1082 (
            .O(N__9112),
            .I(\Lab_UT.scdp.lsBitsD_6 ));
    InMux I__1081 (
            .O(N__9109),
            .I(N__9097));
    InMux I__1080 (
            .O(N__9108),
            .I(N__9097));
    InMux I__1079 (
            .O(N__9107),
            .I(N__9097));
    InMux I__1078 (
            .O(N__9106),
            .I(N__9097));
    LocalMux I__1077 (
            .O(N__9097),
            .I(N__9094));
    Odrv4 I__1076 (
            .O(N__9094),
            .I(\Lab_UT.scdp.d2eData_3_6 ));
    CascadeMux I__1075 (
            .O(N__9091),
            .I(\Lab_UT.scdp.d2eData_3_6_cascade_ ));
    InMux I__1074 (
            .O(N__9088),
            .I(N__9085));
    LocalMux I__1073 (
            .O(N__9085),
            .I(\Lab_UT.scdp.u0.byteToDecrypt_6 ));
    InMux I__1072 (
            .O(N__9082),
            .I(N__9079));
    LocalMux I__1071 (
            .O(N__9079),
            .I(N__9076));
    Span4Mux_v I__1070 (
            .O(N__9076),
            .I(N__9073));
    Odrv4 I__1069 (
            .O(N__9073),
            .I(\ufifo.sb_ram512x8_inst_RNILSN11 ));
    CascadeMux I__1068 (
            .O(N__9070),
            .I(\ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0_cascade_ ));
    InMux I__1067 (
            .O(N__9067),
            .I(N__9060));
    InMux I__1066 (
            .O(N__9066),
            .I(N__9060));
    InMux I__1065 (
            .O(N__9065),
            .I(N__9057));
    LocalMux I__1064 (
            .O(N__9060),
            .I(N__9049));
    LocalMux I__1063 (
            .O(N__9057),
            .I(N__9049));
    InMux I__1062 (
            .O(N__9056),
            .I(N__9044));
    InMux I__1061 (
            .O(N__9055),
            .I(N__9041));
    InMux I__1060 (
            .O(N__9054),
            .I(N__9038));
    Span4Mux_h I__1059 (
            .O(N__9049),
            .I(N__9035));
    InMux I__1058 (
            .O(N__9048),
            .I(N__9030));
    InMux I__1057 (
            .O(N__9047),
            .I(N__9030));
    LocalMux I__1056 (
            .O(N__9044),
            .I(ufifo_utb_txdata_sm0_0));
    LocalMux I__1055 (
            .O(N__9041),
            .I(ufifo_utb_txdata_sm0_0));
    LocalMux I__1054 (
            .O(N__9038),
            .I(ufifo_utb_txdata_sm0_0));
    Odrv4 I__1053 (
            .O(N__9035),
            .I(ufifo_utb_txdata_sm0_0));
    LocalMux I__1052 (
            .O(N__9030),
            .I(ufifo_utb_txdata_sm0_0));
    InMux I__1051 (
            .O(N__9019),
            .I(N__9016));
    LocalMux I__1050 (
            .O(N__9016),
            .I(N__9013));
    Odrv4 I__1049 (
            .O(N__9013),
            .I(utb_txdata_2));
    InMux I__1048 (
            .O(N__9010),
            .I(N__9007));
    LocalMux I__1047 (
            .O(N__9007),
            .I(N__9004));
    Span12Mux_s3_h I__1046 (
            .O(N__9004),
            .I(N__9001));
    Odrv12 I__1045 (
            .O(N__9001),
            .I(\ufifo.txdataDZ0Z_1 ));
    InMux I__1044 (
            .O(N__8998),
            .I(N__8995));
    LocalMux I__1043 (
            .O(N__8995),
            .I(N__8992));
    Odrv4 I__1042 (
            .O(N__8992),
            .I(\Lab_UT.scdp.msBitsi.msBitsD_1 ));
    InMux I__1041 (
            .O(N__8989),
            .I(N__8986));
    LocalMux I__1040 (
            .O(N__8986),
            .I(\Lab_UT.scdp.msBitsi.q_esr_RNI5NL8Z0Z_1 ));
    InMux I__1039 (
            .O(N__8983),
            .I(N__8980));
    LocalMux I__1038 (
            .O(N__8980),
            .I(N__8977));
    Span4Mux_s3_h I__1037 (
            .O(N__8977),
            .I(N__8974));
    Odrv4 I__1036 (
            .O(N__8974),
            .I(\ufifo.txdataDZ0Z_5 ));
    CEMux I__1035 (
            .O(N__8971),
            .I(N__8968));
    LocalMux I__1034 (
            .O(N__8968),
            .I(N__8965));
    Odrv12 I__1033 (
            .O(N__8965),
            .I(\Lab_UT.scdp.u2.sccEldByte_0 ));
    CascadeMux I__1032 (
            .O(N__8962),
            .I(\Lab_UT.scdp.N_52_cascade_ ));
    InMux I__1031 (
            .O(N__8959),
            .I(N__8956));
    LocalMux I__1030 (
            .O(N__8956),
            .I(\Lab_UT.scdp.msBitsi.msBitsDZ0Z_0 ));
    InMux I__1029 (
            .O(N__8953),
            .I(N__8947));
    InMux I__1028 (
            .O(N__8952),
            .I(N__8947));
    LocalMux I__1027 (
            .O(N__8947),
            .I(N__8944));
    Span4Mux_h I__1026 (
            .O(N__8944),
            .I(N__8941));
    Odrv4 I__1025 (
            .O(N__8941),
            .I(\Lab_UT.scdp.byteToEncrypt_4 ));
    CascadeMux I__1024 (
            .O(N__8938),
            .I(N__8935));
    InMux I__1023 (
            .O(N__8935),
            .I(N__8932));
    LocalMux I__1022 (
            .O(N__8932),
            .I(\Lab_UT.scdp.b2a0.N_55 ));
    InMux I__1021 (
            .O(N__8929),
            .I(N__8917));
    InMux I__1020 (
            .O(N__8928),
            .I(N__8917));
    InMux I__1019 (
            .O(N__8927),
            .I(N__8917));
    InMux I__1018 (
            .O(N__8926),
            .I(N__8917));
    LocalMux I__1017 (
            .O(N__8917),
            .I(\Lab_UT.scdp.d2eData_5 ));
    CascadeMux I__1016 (
            .O(N__8914),
            .I(\Lab_UT.scdp.b2a0.N_55_cascade_ ));
    CascadeMux I__1015 (
            .O(N__8911),
            .I(\Lab_UT.scdp.a2b.val_0_0Z0Z_3_cascade_ ));
    InMux I__1014 (
            .O(N__8908),
            .I(N__8905));
    LocalMux I__1013 (
            .O(N__8905),
            .I(N__8902));
    Odrv4 I__1012 (
            .O(N__8902),
            .I(\Lab_UT.scdp.msBitsi.q_esr_RNIF1M8Z0Z_6 ));
    InMux I__1011 (
            .O(N__8899),
            .I(N__8896));
    LocalMux I__1010 (
            .O(N__8896),
            .I(\Lab_UT.scdp.msBitsi.q_esr_RNIQQ8EZ0Z_0 ));
    InMux I__1009 (
            .O(N__8893),
            .I(N__8890));
    LocalMux I__1008 (
            .O(N__8890),
            .I(N__8887));
    Span4Mux_v I__1007 (
            .O(N__8887),
            .I(N__8884));
    Odrv4 I__1006 (
            .O(N__8884),
            .I(\resetGen.escKey_0Z0Z_0 ));
    InMux I__1005 (
            .O(N__8881),
            .I(N__8878));
    LocalMux I__1004 (
            .O(N__8878),
            .I(\Lab_UT.scdp.msBitsi.msBitsD_6 ));
    InMux I__1003 (
            .O(N__8875),
            .I(N__8872));
    LocalMux I__1002 (
            .O(N__8872),
            .I(N__8869));
    Span4Mux_v I__1001 (
            .O(N__8869),
            .I(N__8866));
    Odrv4 I__1000 (
            .O(N__8866),
            .I(\Lab_UT.scdp.u2.byteToEncryptZ0Z_5 ));
    CascadeMux I__999 (
            .O(N__8863),
            .I(\Lab_UT.scdp.d2eData_5_cascade_ ));
    CascadeMux I__998 (
            .O(N__8860),
            .I(N__8856));
    InMux I__997 (
            .O(N__8859),
            .I(N__8845));
    InMux I__996 (
            .O(N__8856),
            .I(N__8845));
    InMux I__995 (
            .O(N__8855),
            .I(N__8845));
    InMux I__994 (
            .O(N__8854),
            .I(N__8845));
    LocalMux I__993 (
            .O(N__8845),
            .I(N__8842));
    Span4Mux_v I__992 (
            .O(N__8842),
            .I(N__8839));
    Odrv4 I__991 (
            .O(N__8839),
            .I(\Lab_UT.scdp.byteToEncrypt_6 ));
    CascadeMux I__990 (
            .O(N__8836),
            .I(\Lab_UT.scdp.q_RNI56C1D_0_cascade_ ));
    InMux I__989 (
            .O(N__8833),
            .I(N__8830));
    LocalMux I__988 (
            .O(N__8830),
            .I(\ufifo.txdataDZ0Z_0 ));
    InMux I__987 (
            .O(N__8827),
            .I(N__8824));
    LocalMux I__986 (
            .O(N__8824),
            .I(N__8821));
    Odrv4 I__985 (
            .O(N__8821),
            .I(\ufifo.txdataDZ0Z_6 ));
    InMux I__984 (
            .O(N__8818),
            .I(N__8813));
    InMux I__983 (
            .O(N__8817),
            .I(N__8808));
    InMux I__982 (
            .O(N__8816),
            .I(N__8808));
    LocalMux I__981 (
            .O(N__8813),
            .I(\resetGen.reset_countZ0Z_2 ));
    LocalMux I__980 (
            .O(N__8808),
            .I(\resetGen.reset_countZ0Z_2 ));
    CascadeMux I__979 (
            .O(N__8803),
            .I(\resetGen.reset_count_2_0_4_cascade_ ));
    InMux I__978 (
            .O(N__8800),
            .I(N__8797));
    LocalMux I__977 (
            .O(N__8797),
            .I(\resetGen.un12_ci ));
    InMux I__976 (
            .O(N__8794),
            .I(N__8791));
    LocalMux I__975 (
            .O(N__8791),
            .I(\resetGen.un23_ci ));
    CascadeMux I__974 (
            .O(N__8788),
            .I(N__8785));
    InMux I__973 (
            .O(N__8785),
            .I(N__8778));
    InMux I__972 (
            .O(N__8784),
            .I(N__8773));
    InMux I__971 (
            .O(N__8783),
            .I(N__8773));
    InMux I__970 (
            .O(N__8782),
            .I(N__8768));
    InMux I__969 (
            .O(N__8781),
            .I(N__8768));
    LocalMux I__968 (
            .O(N__8778),
            .I(N__8763));
    LocalMux I__967 (
            .O(N__8773),
            .I(N__8763));
    LocalMux I__966 (
            .O(N__8768),
            .I(N__8760));
    Span4Mux_h I__965 (
            .O(N__8763),
            .I(N__8757));
    Span4Mux_h I__964 (
            .O(N__8760),
            .I(N__8754));
    Odrv4 I__963 (
            .O(N__8757),
            .I(\resetGen.escKeyZ0 ));
    Odrv4 I__962 (
            .O(N__8754),
            .I(\resetGen.escKeyZ0 ));
    InMux I__961 (
            .O(N__8749),
            .I(N__8743));
    InMux I__960 (
            .O(N__8748),
            .I(N__8743));
    LocalMux I__959 (
            .O(N__8743),
            .I(\resetGen.reset_countZ0Z_3 ));
    InMux I__958 (
            .O(N__8740),
            .I(bfn_4_4_0_));
    CascadeMux I__957 (
            .O(N__8737),
            .I(\resetGen.un12_ci_cascade_ ));
    CascadeMux I__956 (
            .O(N__8734),
            .I(N__8731));
    InMux I__955 (
            .O(N__8731),
            .I(N__8728));
    LocalMux I__954 (
            .O(N__8728),
            .I(N__8724));
    InMux I__953 (
            .O(N__8727),
            .I(N__8720));
    Span4Mux_v I__952 (
            .O(N__8724),
            .I(N__8717));
    InMux I__951 (
            .O(N__8723),
            .I(N__8714));
    LocalMux I__950 (
            .O(N__8720),
            .I(N__8711));
    Odrv4 I__949 (
            .O(N__8717),
            .I(\ufifo.fifo.wraddrZ0Z_6 ));
    LocalMux I__948 (
            .O(N__8714),
            .I(\ufifo.fifo.wraddrZ0Z_6 ));
    Odrv4 I__947 (
            .O(N__8711),
            .I(\ufifo.fifo.wraddrZ0Z_6 ));
    CascadeMux I__946 (
            .O(N__8704),
            .I(N__8701));
    InMux I__945 (
            .O(N__8701),
            .I(N__8698));
    LocalMux I__944 (
            .O(N__8698),
            .I(N__8694));
    InMux I__943 (
            .O(N__8697),
            .I(N__8690));
    Span4Mux_v I__942 (
            .O(N__8694),
            .I(N__8687));
    InMux I__941 (
            .O(N__8693),
            .I(N__8684));
    LocalMux I__940 (
            .O(N__8690),
            .I(N__8681));
    Odrv4 I__939 (
            .O(N__8687),
            .I(\ufifo.fifo.rdaddrZ0Z_7 ));
    LocalMux I__938 (
            .O(N__8684),
            .I(\ufifo.fifo.rdaddrZ0Z_7 ));
    Odrv12 I__937 (
            .O(N__8681),
            .I(\ufifo.fifo.rdaddrZ0Z_7 ));
    CascadeMux I__936 (
            .O(N__8674),
            .I(N__8671));
    InMux I__935 (
            .O(N__8671),
            .I(N__8667));
    CascadeMux I__934 (
            .O(N__8670),
            .I(N__8664));
    LocalMux I__933 (
            .O(N__8667),
            .I(N__8660));
    InMux I__932 (
            .O(N__8664),
            .I(N__8657));
    InMux I__931 (
            .O(N__8663),
            .I(N__8654));
    Span4Mux_v I__930 (
            .O(N__8660),
            .I(N__8649));
    LocalMux I__929 (
            .O(N__8657),
            .I(N__8649));
    LocalMux I__928 (
            .O(N__8654),
            .I(\ufifo.fifo.wraddrZ0Z_7 ));
    Odrv4 I__927 (
            .O(N__8649),
            .I(\ufifo.fifo.wraddrZ0Z_7 ));
    CascadeMux I__926 (
            .O(N__8644),
            .I(N__8641));
    InMux I__925 (
            .O(N__8641),
            .I(N__8638));
    LocalMux I__924 (
            .O(N__8638),
            .I(N__8635));
    Span4Mux_v I__923 (
            .O(N__8635),
            .I(N__8630));
    InMux I__922 (
            .O(N__8634),
            .I(N__8627));
    InMux I__921 (
            .O(N__8633),
            .I(N__8624));
    Sp12to4 I__920 (
            .O(N__8630),
            .I(N__8619));
    LocalMux I__919 (
            .O(N__8627),
            .I(N__8619));
    LocalMux I__918 (
            .O(N__8624),
            .I(\ufifo.fifo.rdaddrZ0Z_6 ));
    Odrv12 I__917 (
            .O(N__8619),
            .I(\ufifo.fifo.rdaddrZ0Z_6 ));
    CascadeMux I__916 (
            .O(N__8614),
            .I(N__8611));
    InMux I__915 (
            .O(N__8611),
            .I(N__8608));
    LocalMux I__914 (
            .O(N__8608),
            .I(N__8603));
    InMux I__913 (
            .O(N__8607),
            .I(N__8600));
    InMux I__912 (
            .O(N__8606),
            .I(N__8597));
    Span4Mux_v I__911 (
            .O(N__8603),
            .I(N__8592));
    LocalMux I__910 (
            .O(N__8600),
            .I(N__8592));
    LocalMux I__909 (
            .O(N__8597),
            .I(\ufifo.fifo.wraddrZ0Z_0 ));
    Odrv4 I__908 (
            .O(N__8592),
            .I(\ufifo.fifo.wraddrZ0Z_0 ));
    CascadeMux I__907 (
            .O(N__8587),
            .I(N__8584));
    InMux I__906 (
            .O(N__8584),
            .I(N__8581));
    LocalMux I__905 (
            .O(N__8581),
            .I(N__8576));
    InMux I__904 (
            .O(N__8580),
            .I(N__8573));
    InMux I__903 (
            .O(N__8579),
            .I(N__8570));
    Sp12to4 I__902 (
            .O(N__8576),
            .I(N__8565));
    LocalMux I__901 (
            .O(N__8573),
            .I(N__8565));
    LocalMux I__900 (
            .O(N__8570),
            .I(\ufifo.fifo.rdaddrZ0Z_8 ));
    Odrv12 I__899 (
            .O(N__8565),
            .I(\ufifo.fifo.rdaddrZ0Z_8 ));
    CascadeMux I__898 (
            .O(N__8560),
            .I(N__8557));
    InMux I__897 (
            .O(N__8557),
            .I(N__8552));
    CascadeMux I__896 (
            .O(N__8556),
            .I(N__8549));
    InMux I__895 (
            .O(N__8555),
            .I(N__8546));
    LocalMux I__894 (
            .O(N__8552),
            .I(N__8543));
    InMux I__893 (
            .O(N__8549),
            .I(N__8540));
    LocalMux I__892 (
            .O(N__8546),
            .I(N__8535));
    Span4Mux_v I__891 (
            .O(N__8543),
            .I(N__8535));
    LocalMux I__890 (
            .O(N__8540),
            .I(N__8532));
    Odrv4 I__889 (
            .O(N__8535),
            .I(\ufifo.fifo.wraddrZ0Z_8 ));
    Odrv4 I__888 (
            .O(N__8532),
            .I(\ufifo.fifo.wraddrZ0Z_8 ));
    CascadeMux I__887 (
            .O(N__8527),
            .I(N__8524));
    InMux I__886 (
            .O(N__8524),
            .I(N__8521));
    LocalMux I__885 (
            .O(N__8521),
            .I(N__8518));
    Span4Mux_v I__884 (
            .O(N__8518),
            .I(N__8513));
    InMux I__883 (
            .O(N__8517),
            .I(N__8510));
    InMux I__882 (
            .O(N__8516),
            .I(N__8507));
    Sp12to4 I__881 (
            .O(N__8513),
            .I(N__8502));
    LocalMux I__880 (
            .O(N__8510),
            .I(N__8502));
    LocalMux I__879 (
            .O(N__8507),
            .I(\ufifo.fifo.rdaddrZ0Z_0 ));
    Odrv12 I__878 (
            .O(N__8502),
            .I(\ufifo.fifo.rdaddrZ0Z_0 ));
    InMux I__877 (
            .O(N__8497),
            .I(N__8485));
    InMux I__876 (
            .O(N__8496),
            .I(N__8485));
    InMux I__875 (
            .O(N__8495),
            .I(N__8485));
    InMux I__874 (
            .O(N__8494),
            .I(N__8485));
    LocalMux I__873 (
            .O(N__8485),
            .I(\resetGen.reset_countZ0Z_0 ));
    InMux I__872 (
            .O(N__8482),
            .I(N__8473));
    InMux I__871 (
            .O(N__8481),
            .I(N__8473));
    InMux I__870 (
            .O(N__8480),
            .I(N__8473));
    LocalMux I__869 (
            .O(N__8473),
            .I(\resetGen.reset_countZ0Z_1 ));
    InMux I__868 (
            .O(N__8470),
            .I(bfn_4_2_0_));
    InMux I__867 (
            .O(N__8467),
            .I(\ufifo.fifo.un1_wraddr_cry_0 ));
    InMux I__866 (
            .O(N__8464),
            .I(\ufifo.fifo.un1_wraddr_cry_1 ));
    InMux I__865 (
            .O(N__8461),
            .I(\ufifo.fifo.un1_wraddr_cry_2 ));
    InMux I__864 (
            .O(N__8458),
            .I(\ufifo.fifo.un1_wraddr_cry_3 ));
    InMux I__863 (
            .O(N__8455),
            .I(\ufifo.fifo.un1_wraddr_cry_4 ));
    InMux I__862 (
            .O(N__8452),
            .I(\ufifo.fifo.un1_wraddr_cry_5 ));
    InMux I__861 (
            .O(N__8449),
            .I(\ufifo.fifo.un1_wraddr_cry_6 ));
    InMux I__860 (
            .O(N__8446),
            .I(N__8443));
    LocalMux I__859 (
            .O(N__8443),
            .I(\Lab_UT.scdp.u2.byteToEncrypt_0 ));
    InMux I__858 (
            .O(N__8440),
            .I(\ufifo.fifo.un1_rdaddr_cry_0 ));
    InMux I__857 (
            .O(N__8437),
            .I(\ufifo.fifo.un1_rdaddr_cry_1 ));
    InMux I__856 (
            .O(N__8434),
            .I(\ufifo.fifo.un1_rdaddr_cry_2 ));
    InMux I__855 (
            .O(N__8431),
            .I(\ufifo.fifo.un1_rdaddr_cry_3 ));
    InMux I__854 (
            .O(N__8428),
            .I(\ufifo.fifo.un1_rdaddr_cry_4 ));
    InMux I__853 (
            .O(N__8425),
            .I(\ufifo.fifo.un1_rdaddr_cry_5 ));
    InMux I__852 (
            .O(N__8422),
            .I(\ufifo.fifo.un1_rdaddr_cry_6 ));
    InMux I__851 (
            .O(N__8419),
            .I(N__8416));
    LocalMux I__850 (
            .O(N__8416),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__849 (
            .O(N__8413),
            .I(N__8410));
    LocalMux I__848 (
            .O(N__8410),
            .I(N__8407));
    Odrv4 I__847 (
            .O(N__8407),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__846 (
            .O(N__8404),
            .I(N__8401));
    LocalMux I__845 (
            .O(N__8401),
            .I(N__8398));
    Odrv4 I__844 (
            .O(N__8398),
            .I(ufifo_utb_txdata_m0_4));
    CascadeMux I__843 (
            .O(N__8395),
            .I(N__8392));
    InMux I__842 (
            .O(N__8392),
            .I(N__8389));
    LocalMux I__841 (
            .O(N__8389),
            .I(N__8386));
    Odrv4 I__840 (
            .O(N__8386),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    CascadeMux I__839 (
            .O(N__8383),
            .I(N__8380));
    InMux I__838 (
            .O(N__8380),
            .I(N__8377));
    LocalMux I__837 (
            .O(N__8377),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    CEMux I__836 (
            .O(N__8374),
            .I(N__8368));
    CEMux I__835 (
            .O(N__8373),
            .I(N__8365));
    CEMux I__834 (
            .O(N__8372),
            .I(N__8362));
    CEMux I__833 (
            .O(N__8371),
            .I(N__8359));
    LocalMux I__832 (
            .O(N__8368),
            .I(N__8354));
    LocalMux I__831 (
            .O(N__8365),
            .I(N__8354));
    LocalMux I__830 (
            .O(N__8362),
            .I(N__8351));
    LocalMux I__829 (
            .O(N__8359),
            .I(N__8348));
    Odrv4 I__828 (
            .O(N__8354),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__827 (
            .O(N__8351),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__826 (
            .O(N__8348),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    CascadeMux I__825 (
            .O(N__8341),
            .I(N__8338));
    InMux I__824 (
            .O(N__8338),
            .I(N__8335));
    LocalMux I__823 (
            .O(N__8335),
            .I(N__8332));
    Odrv4 I__822 (
            .O(N__8332),
            .I(\Lab_UT.scdp.byteToEncrypt_7 ));
    CascadeMux I__821 (
            .O(N__8329),
            .I(\ufifo.un4_rxDataValidNoEscZ0Z_1_cascade_ ));
    InMux I__820 (
            .O(N__8326),
            .I(N__8323));
    LocalMux I__819 (
            .O(N__8323),
            .I(\ufifo.rxDataValidNoEscZ0 ));
    CascadeMux I__818 (
            .O(N__8320),
            .I(N__8317));
    InMux I__817 (
            .O(N__8317),
            .I(N__8314));
    LocalMux I__816 (
            .O(N__8314),
            .I(N__8311));
    Odrv4 I__815 (
            .O(N__8311),
            .I(\ufifo.fifo.fifo_txdata_3 ));
    InMux I__814 (
            .O(N__8308),
            .I(N__8305));
    LocalMux I__813 (
            .O(N__8305),
            .I(\ufifo.fifo.fifo_txdata_4 ));
    CascadeMux I__812 (
            .O(N__8302),
            .I(N__8299));
    InMux I__811 (
            .O(N__8299),
            .I(N__8296));
    LocalMux I__810 (
            .O(N__8296),
            .I(N__8293));
    Odrv4 I__809 (
            .O(N__8293),
            .I(\ufifo.utb_txdata_m0_0 ));
    InMux I__808 (
            .O(N__8290),
            .I(N__8287));
    LocalMux I__807 (
            .O(N__8287),
            .I(utb_txdata_0));
    CascadeMux I__806 (
            .O(N__8284),
            .I(N__8281));
    InMux I__805 (
            .O(N__8281),
            .I(N__8275));
    InMux I__804 (
            .O(N__8280),
            .I(N__8275));
    LocalMux I__803 (
            .O(N__8275),
            .I(Lab_UT_dk_de_cr_2_reti));
    InMux I__802 (
            .O(N__8272),
            .I(N__8269));
    LocalMux I__801 (
            .O(N__8269),
            .I(ufifo_utb_txdata_m0_3));
    CascadeMux I__800 (
            .O(N__8266),
            .I(\ufifo.sb_ram512x8_inst_RNIKRN11_cascade_ ));
    InMux I__799 (
            .O(N__8263),
            .I(N__8260));
    LocalMux I__798 (
            .O(N__8260),
            .I(\ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0 ));
    InMux I__797 (
            .O(N__8257),
            .I(N__8254));
    LocalMux I__796 (
            .O(N__8254),
            .I(utb_txdata_1));
    InMux I__795 (
            .O(N__8251),
            .I(N__8248));
    LocalMux I__794 (
            .O(N__8248),
            .I(\ufifo.fifo.fifo_txdata_0 ));
    InMux I__793 (
            .O(N__8245),
            .I(N__8242));
    LocalMux I__792 (
            .O(N__8242),
            .I(N__8239));
    Odrv4 I__791 (
            .O(N__8239),
            .I(\ufifo.fifo.fifo_txdata_6 ));
    InMux I__790 (
            .O(N__8236),
            .I(N__8233));
    LocalMux I__789 (
            .O(N__8233),
            .I(N__8230));
    Odrv4 I__788 (
            .O(N__8230),
            .I(\ufifo.fifo.fifo_txdata_5 ));
    InMux I__787 (
            .O(N__8227),
            .I(N__8224));
    LocalMux I__786 (
            .O(N__8224),
            .I(ufifo_utb_txdata_m0_5));
    InMux I__785 (
            .O(N__8221),
            .I(N__8218));
    LocalMux I__784 (
            .O(N__8218),
            .I(\ufifo.fifo.fifo_txdata_7 ));
    InMux I__783 (
            .O(N__8215),
            .I(N__8212));
    LocalMux I__782 (
            .O(N__8212),
            .I(ufifo_utb_txdata_m0_7));
    InMux I__781 (
            .O(N__8209),
            .I(N__8206));
    LocalMux I__780 (
            .O(N__8206),
            .I(ufifo_utb_txdata_m0_6));
    CascadeMux I__779 (
            .O(N__8203),
            .I(N__8200));
    InMux I__778 (
            .O(N__8200),
            .I(N__8197));
    LocalMux I__777 (
            .O(N__8197),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CascadeMux I__776 (
            .O(N__8194),
            .I(N__8191));
    InMux I__775 (
            .O(N__8191),
            .I(N__8188));
    LocalMux I__774 (
            .O(N__8188),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__773 (
            .O(N__8185),
            .I(N__8182));
    LocalMux I__772 (
            .O(N__8182),
            .I(\buart.Z_tx.counter_RNIVE1P1_1 ));
    InMux I__771 (
            .O(N__8179),
            .I(\buart.Z_tx.un1_bitcount_cry_0 ));
    InMux I__770 (
            .O(N__8176),
            .I(N__8173));
    LocalMux I__769 (
            .O(N__8173),
            .I(\buart.Z_tx.counter_RNIVE1P1_0_1 ));
    InMux I__768 (
            .O(N__8170),
            .I(\buart.Z_tx.un1_bitcount_cry_1 ));
    InMux I__767 (
            .O(N__8167),
            .I(N__8164));
    LocalMux I__766 (
            .O(N__8164),
            .I(\buart.Z_tx.un1_bitcount_axb_3 ));
    InMux I__765 (
            .O(N__8161),
            .I(\buart.Z_tx.un1_bitcount_cry_2 ));
    CascadeMux I__764 (
            .O(N__8158),
            .I(N__8155));
    InMux I__763 (
            .O(N__8155),
            .I(N__8152));
    LocalMux I__762 (
            .O(N__8152),
            .I(\buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0 ));
    CascadeMux I__761 (
            .O(N__8149),
            .I(N__8146));
    InMux I__760 (
            .O(N__8146),
            .I(N__8143));
    LocalMux I__759 (
            .O(N__8143),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    InMux I__758 (
            .O(N__8140),
            .I(N__8135));
    InMux I__757 (
            .O(N__8139),
            .I(N__8130));
    InMux I__756 (
            .O(N__8138),
            .I(N__8130));
    LocalMux I__755 (
            .O(N__8135),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__754 (
            .O(N__8130),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    InMux I__753 (
            .O(N__8125),
            .I(N__8122));
    LocalMux I__752 (
            .O(N__8122),
            .I(\ufifo.fifo.fifo_txdata_2 ));
    InMux I__751 (
            .O(N__8119),
            .I(N__8116));
    LocalMux I__750 (
            .O(N__8116),
            .I(\ufifo.fifo.fifo_txdata_1 ));
    InMux I__749 (
            .O(N__8113),
            .I(N__8110));
    LocalMux I__748 (
            .O(N__8110),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__747 (
            .O(N__8107),
            .I(N__8104));
    LocalMux I__746 (
            .O(N__8104),
            .I(N__8101));
    IoSpan4Mux I__745 (
            .O(N__8101),
            .I(N__8098));
    Odrv4 I__744 (
            .O(N__8098),
            .I(o_serial_data_c));
    InMux I__743 (
            .O(N__8095),
            .I(N__8092));
    LocalMux I__742 (
            .O(N__8092),
            .I(uart_RXD));
    InMux I__741 (
            .O(N__8089),
            .I(N__8083));
    InMux I__740 (
            .O(N__8088),
            .I(N__8083));
    LocalMux I__739 (
            .O(N__8083),
            .I(N__8080));
    Odrv4 I__738 (
            .O(N__8080),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    InMux I__737 (
            .O(N__8077),
            .I(N__8074));
    LocalMux I__736 (
            .O(N__8074),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3 ));
    CascadeMux I__735 (
            .O(N__8071),
            .I(N__8067));
    InMux I__734 (
            .O(N__8070),
            .I(N__8059));
    InMux I__733 (
            .O(N__8067),
            .I(N__8059));
    InMux I__732 (
            .O(N__8066),
            .I(N__8059));
    LocalMux I__731 (
            .O(N__8059),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    IoInMux I__730 (
            .O(N__8056),
            .I(N__8053));
    LocalMux I__729 (
            .O(N__8053),
            .I(N__8050));
    IoSpan4Mux I__728 (
            .O(N__8050),
            .I(N__8047));
    Span4Mux_s0_h I__727 (
            .O(N__8047),
            .I(N__8044));
    Odrv4 I__726 (
            .O(N__8044),
            .I(\buart.Z_rx.N_41_i ));
    InMux I__725 (
            .O(N__8041),
            .I(N__8035));
    InMux I__724 (
            .O(N__8040),
            .I(N__8032));
    InMux I__723 (
            .O(N__8039),
            .I(N__8027));
    InMux I__722 (
            .O(N__8038),
            .I(N__8027));
    LocalMux I__721 (
            .O(N__8035),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__720 (
            .O(N__8032),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__719 (
            .O(N__8027),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__718 (
            .O(N__8020),
            .I(N__8017));
    LocalMux I__717 (
            .O(N__8017),
            .I(N__8014));
    Odrv4 I__716 (
            .O(N__8014),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    CascadeMux I__715 (
            .O(N__8011),
            .I(N__8006));
    InMux I__714 (
            .O(N__8010),
            .I(N__8003));
    InMux I__713 (
            .O(N__8009),
            .I(N__8000));
    InMux I__712 (
            .O(N__8006),
            .I(N__7997));
    LocalMux I__711 (
            .O(N__8003),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__710 (
            .O(N__8000),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__709 (
            .O(N__7997),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    InMux I__708 (
            .O(N__7990),
            .I(N__7987));
    LocalMux I__707 (
            .O(N__7987),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__706 (
            .O(N__7984),
            .I(N__7981));
    LocalMux I__705 (
            .O(N__7981),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    CascadeMux I__704 (
            .O(N__7978),
            .I(N__7975));
    InMux I__703 (
            .O(N__7975),
            .I(N__7970));
    InMux I__702 (
            .O(N__7974),
            .I(N__7965));
    InMux I__701 (
            .O(N__7973),
            .I(N__7965));
    LocalMux I__700 (
            .O(N__7970),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__699 (
            .O(N__7965),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    InMux I__698 (
            .O(N__7960),
            .I(N__7954));
    InMux I__697 (
            .O(N__7959),
            .I(N__7947));
    InMux I__696 (
            .O(N__7958),
            .I(N__7947));
    InMux I__695 (
            .O(N__7957),
            .I(N__7947));
    LocalMux I__694 (
            .O(N__7954),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__693 (
            .O(N__7947),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__692 (
            .O(N__7942),
            .I(N__7938));
    InMux I__691 (
            .O(N__7941),
            .I(N__7935));
    InMux I__690 (
            .O(N__7938),
            .I(N__7932));
    LocalMux I__689 (
            .O(N__7935),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__688 (
            .O(N__7932),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    InMux I__687 (
            .O(N__7927),
            .I(N__7924));
    LocalMux I__686 (
            .O(N__7924),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    InMux I__685 (
            .O(N__7921),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__684 (
            .O(N__7918),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__683 (
            .O(N__7915),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    InMux I__682 (
            .O(N__7912),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    InMux I__681 (
            .O(N__7909),
            .I(N__7903));
    InMux I__680 (
            .O(N__7908),
            .I(N__7903));
    LocalMux I__679 (
            .O(N__7903),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    InMux I__678 (
            .O(N__7900),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__677 (
            .O(N__7897),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__676 (
            .O(N__7894),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__675 (
            .O(N__7891),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__674 (
            .O(N__7888),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    InMux I__673 (
            .O(N__7885),
            .I(N__7879));
    InMux I__672 (
            .O(N__7884),
            .I(N__7879));
    LocalMux I__671 (
            .O(N__7879),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__670 (
            .O(N__7876),
            .I(N__7873));
    InMux I__669 (
            .O(N__7873),
            .I(N__7867));
    InMux I__668 (
            .O(N__7872),
            .I(N__7867));
    LocalMux I__667 (
            .O(N__7867),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    CascadeMux I__666 (
            .O(N__7864),
            .I(N__7860));
    CascadeMux I__665 (
            .O(N__7863),
            .I(N__7857));
    InMux I__664 (
            .O(N__7860),
            .I(N__7852));
    InMux I__663 (
            .O(N__7857),
            .I(N__7852));
    LocalMux I__662 (
            .O(N__7852),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    InMux I__661 (
            .O(N__7849),
            .I(N__7843));
    InMux I__660 (
            .O(N__7848),
            .I(N__7843));
    LocalMux I__659 (
            .O(N__7843),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    IoInMux I__658 (
            .O(N__7840),
            .I(N__7837));
    LocalMux I__657 (
            .O(N__7837),
            .I(N__7834));
    Span12Mux_s1_v I__656 (
            .O(N__7834),
            .I(N__7831));
    Span12Mux_v I__655 (
            .O(N__7831),
            .I(N__7828));
    Odrv12 I__654 (
            .O(N__7828),
            .I(\latticehx1k_pll_inst.clk ));
    IoInMux I__653 (
            .O(N__7825),
            .I(N__7822));
    LocalMux I__652 (
            .O(N__7822),
            .I(N__7819));
    IoSpan4Mux I__651 (
            .O(N__7819),
            .I(N__7816));
    Odrv4 I__650 (
            .O(N__7816),
            .I(clk_in_c));
    defparam IN_MUX_bfv_2_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_5_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_4_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_3_0_));
    defparam IN_MUX_bfv_4_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_4_0_ (
            .carryinitin(\ufifo.fifo.un1_wraddr_cry_7 ),
            .carryinitout(bfn_4_4_0_));
    defparam IN_MUX_bfv_4_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_1_0_));
    defparam IN_MUX_bfv_4_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_2_0_ (
            .carryinitin(\ufifo.fifo.un1_rdaddr_cry_7 ),
            .carryinitout(bfn_4_2_0_));
    ICE_GB \buart.Z_rx.bitcount_es_RNIV4M42_0_4  (
            .USERSIGNALTOGLOBALBUFFER(N__8056),
            .GLOBALBUFFEROUTPUT(N_41_i_g));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__7840),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__12676),
            .GLOBALBUFFEROUTPUT(\Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_g ));
    ICE_GB \resetGen.rst_0_iso_RNITVH4  (
            .USERSIGNALTOGLOBALBUFFER(N__14086),
            .GLOBALBUFFEROUTPUT(resetGen_rst_0_iso_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_3_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_3_0  (
            .in0(_gnd_net_),
            .in1(N__7960),
            .in2(N__7978),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_3_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_3_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_1_3_1  (
            .in0(_gnd_net_),
            .in1(N__7849),
            .in2(_gnd_net_),
            .in3(N__7900),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__22699),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_3_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_3_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_3_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_1_3_2  (
            .in0(N__12094),
            .in1(_gnd_net_),
            .in2(N__7876),
            .in3(N__7897),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__22699),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_3_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_3_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(N__7941),
            .in2(_gnd_net_),
            .in3(N__7894),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__22699),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_3_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_3_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_1_3_4  (
            .in0(N__12095),
            .in1(N__7885),
            .in2(_gnd_net_),
            .in3(N__7891),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__22699),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_3_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_3_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_3_5 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_1_3_5  (
            .in0(_gnd_net_),
            .in1(N__12093),
            .in2(N__7864),
            .in3(N__7888),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22699),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIGU38_6_LC_1_3_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIGU38_6_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIGU38_6_LC_1_3_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIGU38_6_LC_1_3_7  (
            .in0(N__7884),
            .in1(N__7872),
            .in2(N__7863),
            .in3(N__7848),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_4_0 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_4_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_4_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_1_4_0  (
            .in0(N__7959),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7974),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22696),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_4_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_4_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_4_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_1_4_6  (
            .in0(N__7958),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22696),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_4_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_4_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_4_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_4_7  (
            .in0(N__7973),
            .in1(N__7957),
            .in2(N__7942),
            .in3(N__7927),
            .lcout(\buart.Z_tx.N_255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1_0_LC_1_5_6 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1_0_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1_0_LC_1_5_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1_0_LC_1_5_6  (
            .in0(N__11374),
            .in1(N__9917),
            .in2(_gnd_net_),
            .in3(N__11462),
            .lcout(\ufifo.crlfdone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_0_LC_1_5_7 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_0_LC_1_5_7 .SEQ_MODE=4'b1000;
    defparam \ufifo.emitcrlf_fsm.cstate_0_LC_1_5_7 .LUT_INIT=16'b0111100000000000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_0_LC_1_5_7  (
            .in0(N__11463),
            .in1(N__11375),
            .in2(N__9931),
            .in3(N__20243),
            .lcout(\ufifo.emitcrlf_fsm.cstateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22693),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_1_6_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_1_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__8039),
            .in2(N__8071),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_1_6_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_1_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__8139),
            .in2(_gnd_net_),
            .in3(N__7921),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_1_6_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_1_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_1_6_2  (
            .in0(N__10367),
            .in1(N__7909),
            .in2(_gnd_net_),
            .in3(N__7918),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__22689),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_1_6_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_1_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(N__8009),
            .in2(_gnd_net_),
            .in3(N__7915),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_1_6_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_1_6_4 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_1_6_4  (
            .in0(N__8089),
            .in1(N__10366),
            .in2(N__10182),
            .in3(N__7912),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22689),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_1_6_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_1_6_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_1_6_5  (
            .in0(N__7908),
            .in1(N__8138),
            .in2(N__8011),
            .in3(N__8066),
            .lcout(\buart.Z_rx.Z_baudgen.ser_clk_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_1_6_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_1_6_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_1_6_6  (
            .in0(N__8088),
            .in1(N__8038),
            .in2(_gnd_net_),
            .in3(N__8077),
            .lcout(\buart.Z_rx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_1_6_7 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_1_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_1_6_7  (
            .in0(N__10365),
            .in1(N__8041),
            .in2(_gnd_net_),
            .in3(N__8070),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22689),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_4_LC_1_7_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_4_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_4_LC_1_7_3 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIV4M42_4_LC_1_7_3  (
            .in0(N__10170),
            .in1(N__10497),
            .in2(N__10408),
            .in3(N__10609),
            .lcout(\buart.Z_rx.N_41_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_1_7_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_1_7_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_1_7_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(N__8040),
            .in2(_gnd_net_),
            .in3(N__10377),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22682),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_1_7_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_1_7_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_1_7_5 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_1_7_5  (
            .in0(N__10171),
            .in1(N__8020),
            .in2(N__10378),
            .in3(N__8010),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22682),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_0_LC_1_7_7 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_0_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_0_LC_1_7_7 .LUT_INIT=16'b1001100111111111;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_0_LC_1_7_7  (
            .in0(N__11386),
            .in1(N__9924),
            .in2(_gnd_net_),
            .in3(N__11467),
            .lcout(ufifo_utb_txdata_sm0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_1_8_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_1_8_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_1_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \buart.Z_tx.shifter_1_LC_1_8_4  (
            .in0(N__7990),
            .in1(N__8290),
            .in2(_gnd_net_),
            .in3(N__12038),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22676),
            .ce(N__8374),
            .sr(N__18063));
    defparam \buart.Z_tx.shifter_6_LC_1_8_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_1_8_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_1_8_6 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \buart.Z_tx.shifter_6_LC_1_8_6  (
            .in0(N__8227),
            .in1(N__9055),
            .in2(N__8194),
            .in3(N__12039),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22676),
            .ce(N__8374),
            .sr(N__18063));
    defparam \buart.Z_tx.shifter_2_LC_1_8_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_1_8_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_1_8_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \buart.Z_tx.shifter_2_LC_1_8_7  (
            .in0(N__12037),
            .in1(N__8413),
            .in2(_gnd_net_),
            .in3(N__8257),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22676),
            .ce(N__8374),
            .sr(N__18063));
    defparam \buart.Z_tx.shifter_0_LC_1_9_2 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_1_9_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_1_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_tx.shifter_0_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__7984),
            .in2(_gnd_net_),
            .in3(N__12051),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22668),
            .ce(N__8371),
            .sr(N__18065));
    defparam \buart.Z_tx.uart_tx_LC_1_9_5 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_1_9_5 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_1_9_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \buart.Z_tx.uart_tx_LC_1_9_5  (
            .in0(N__12050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8113),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22668),
            .ce(N__8371),
            .sr(N__18065));
    defparam \buart.Z_rx.hh_1_LC_1_10_6 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_1_10_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_1_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10212),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22664),
            .ce(),
            .sr(N__18066));
    defparam \buart.Z_rx.hh_0_LC_1_11_7 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_1_11_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8095),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22655),
            .ce(),
            .sr(N__18067));
    defparam \ufifo.tx_fsm.cstate_3_LC_2_3_1 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_3_LC_2_3_1 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_3_LC_2_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ufifo.tx_fsm.cstate_3_LC_2_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10024),
            .lcout(\ufifo.tx_fsm.fifo_txdata_rdy ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22697),
            .ce(),
            .sr(N__9959));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_1_LC_2_4_2 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_1_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_1_LC_2_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_1_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(N__12086),
            .in2(_gnd_net_),
            .in3(N__12176),
            .lcout(\buart.Z_tx.counter_RNIVE1P1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_0_1_LC_2_4_3 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_0_1_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_0_1_LC_2_4_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_0_1_LC_2_4_3  (
            .in0(N__12177),
            .in1(_gnd_net_),
            .in2(N__12103),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.counter_RNIVE1P1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.state_ret_5_RNIAFUE_LC_2_4_4 .C_ON=1'b0;
    defparam \resetGen.state_ret_5_RNIAFUE_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \resetGen.state_ret_5_RNIAFUE_LC_2_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.state_ret_5_RNIAFUE_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20271),
            .lcout(rst_i_3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_2_4_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_2_4_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_2_4_7  (
            .in0(N__12178),
            .in1(_gnd_net_),
            .in2(N__12104),
            .in3(N__10095),
            .lcout(\buart.Z_tx.un1_bitcount_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_LC_2_5_0 .C_ON=1'b1;
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_LC_2_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.un1_bitcount_cry_0_0_c_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(N__11968),
            .in2(N__8158),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_5_0_),
            .carryout(\buart.Z_tx.un1_bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_1_LC_2_5_1 .C_ON=1'b1;
    defparam \buart.Z_tx.bitcount_1_LC_2_5_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_2_5_1 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_2_5_1  (
            .in0(N__12048),
            .in1(N__8185),
            .in2(N__10117),
            .in3(N__8179),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(\buart.Z_tx.un1_bitcount_cry_0 ),
            .carryout(\buart.Z_tx.un1_bitcount_cry_1 ),
            .clk(N__22690),
            .ce(),
            .sr(N__18070));
    defparam \buart.Z_tx.bitcount_2_LC_2_5_2 .C_ON=1'b1;
    defparam \buart.Z_tx.bitcount_2_LC_2_5_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_2_5_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_2_5_2  (
            .in0(N__12047),
            .in1(N__8176),
            .in2(N__10135),
            .in3(N__8170),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.un1_bitcount_cry_1 ),
            .carryout(\buart.Z_tx.un1_bitcount_cry_2 ),
            .clk(N__22690),
            .ce(),
            .sr(N__18070));
    defparam \buart.Z_tx.bitcount_3_LC_2_5_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_2_5_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_2_5_3 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_2_5_3  (
            .in0(N__12049),
            .in1(N__8167),
            .in2(_gnd_net_),
            .in3(N__8161),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22690),
            .ce(),
            .sr(N__18070));
    defparam \resetGen.rst_0_iso_LC_2_6_0 .C_ON=1'b0;
    defparam \resetGen.rst_0_iso_LC_2_6_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_0_iso_LC_2_6_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \resetGen.rst_0_iso_LC_2_6_0  (
            .in0(N__22761),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(resetGen_rst_0_iso),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22683),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_RNO_LC_2_6_3 .C_ON=1'b0;
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_RNO_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_RNO_LC_2_6_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \buart.Z_tx.un1_bitcount_cry_0_0_c_RNO_LC_2_6_3  (
            .in0(N__12096),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12158),
            .lcout(\buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_6_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_6_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_6_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_2_6_4  (
            .in0(N__10364),
            .in1(N__8140),
            .in2(N__8149),
            .in3(N__10178),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22683),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_LC_2_6_5 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_LC_2_6_5 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_LC_2_6_5  (
            .in0(N__11387),
            .in1(N__9916),
            .in2(_gnd_net_),
            .in3(N__11469),
            .lcout(\ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNILSN11_LC_2_6_7 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNILSN11_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNILSN11_LC_2_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNILSN11_LC_2_6_7  (
            .in0(N__11242),
            .in1(N__8125),
            .in2(_gnd_net_),
            .in3(N__15686),
            .lcout(\ufifo.sb_ram512x8_inst_RNILSN11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIKRN11_LC_2_7_0 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIKRN11_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIKRN11_LC_2_7_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNIKRN11_LC_2_7_0  (
            .in0(N__15771),
            .in1(N__11262),
            .in2(_gnd_net_),
            .in3(N__8119),
            .lcout(),
            .ltout(\ufifo.sb_ram512x8_inst_RNIKRN11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIQ6FP3_0_LC_2_7_1 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIQ6FP3_0_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIQ6FP3_0_LC_2_7_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIQ6FP3_0_LC_2_7_1  (
            .in0(N__9048),
            .in1(_gnd_net_),
            .in2(N__8266),
            .in3(N__8263),
            .lcout(utb_txdata_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIJQN11_LC_2_7_2 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIJQN11_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIJQN11_LC_2_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNIJQN11_LC_2_7_2  (
            .in0(N__11263),
            .in1(N__8251),
            .in2(_gnd_net_),
            .in3(N__16166),
            .lcout(\ufifo.utb_txdata_m0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIP0O11_LC_2_7_3 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIP0O11_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIP0O11_LC_2_7_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNIP0O11_LC_2_7_3  (
            .in0(N__8245),
            .in1(N__11267),
            .in2(_gnd_net_),
            .in3(N__17074),
            .lcout(ufifo_utb_txdata_m0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNIA4BA7_3_LC_2_7_4 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNIA4BA7_3_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNIA4BA7_3_LC_2_7_4 .LUT_INIT=16'b0000000010001100;
    LogicCell40 \ufifo.tx_fsm.cstate_RNIA4BA7_3_LC_2_7_4  (
            .in0(N__11264),
            .in1(N__9047),
            .in2(N__9510),
            .in3(N__8326),
            .lcout(ufifo_utb_txdata_rdy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIOVN11_LC_2_7_5 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIOVN11_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIOVN11_LC_2_7_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNIOVN11_LC_2_7_5  (
            .in0(N__8236),
            .in1(N__11266),
            .in2(_gnd_net_),
            .in3(N__13437),
            .lcout(ufifo_utb_txdata_m0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIQ1O11_LC_2_7_7 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIQ1O11_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIQ1O11_LC_2_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNIQ1O11_LC_2_7_7  (
            .in0(N__8221),
            .in1(N__11265),
            .in2(_gnd_net_),
            .in3(N__16964),
            .lcout(ufifo_utb_txdata_m0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_8_LC_2_8_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_2_8_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_2_8_1 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \buart.Z_tx.shifter_8_LC_2_8_1  (
            .in0(N__8215),
            .in1(N__9054),
            .in2(_gnd_net_),
            .in3(N__12036),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22669),
            .ce(N__8373),
            .sr(N__18064));
    defparam \buart.Z_tx.shifter_7_LC_2_8_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_2_8_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_2_8_4 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \buart.Z_tx.shifter_7_LC_2_8_4  (
            .in0(N__12035),
            .in1(N__8209),
            .in2(N__8203),
            .in3(N__9056),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22669),
            .ce(N__8373),
            .sr(N__18064));
    defparam \ufifo.un4_rxDataValidNoEsc_1_LC_2_8_5 .C_ON=1'b0;
    defparam \ufifo.un4_rxDataValidNoEsc_1_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \ufifo.un4_rxDataValidNoEsc_1_LC_2_8_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \ufifo.un4_rxDataValidNoEsc_1_LC_2_8_5  (
            .in0(N__13318),
            .in1(N__16955),
            .in2(N__15702),
            .in3(N__11680),
            .lcout(),
            .ltout(\ufifo.un4_rxDataValidNoEscZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.rxDataValidNoEsc_LC_2_8_6 .C_ON=1'b0;
    defparam \ufifo.rxDataValidNoEsc_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \ufifo.rxDataValidNoEsc_LC_2_8_6 .LUT_INIT=16'b1011111100000000;
    LogicCell40 \ufifo.rxDataValidNoEsc_LC_2_8_6  (
            .in0(N__11592),
            .in1(N__8280),
            .in2(N__8329),
            .in3(N__20809),
            .lcout(\ufifo.rxDataValidNoEscZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_LC_2_8_7 .C_ON=1'b0;
    defparam \resetGen.escKey_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_LC_2_8_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \resetGen.escKey_LC_2_8_7  (
            .in0(N__20810),
            .in1(N__8893),
            .in2(N__8284),
            .in3(N__11593),
            .lcout(\resetGen.escKeyZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_3_LC_2_9_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_3_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_3_LC_2_9_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_3_LC_2_9_0  (
            .in0(N__11041),
            .in1(N__10798),
            .in2(N__8341),
            .in3(N__10954),
            .lcout(\Lab_UT.scdp.N_48_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIMTN11_LC_2_9_1 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIMTN11_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIMTN11_LC_2_9_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNIMTN11_LC_2_9_1  (
            .in0(N__11922),
            .in1(_gnd_net_),
            .in2(N__8320),
            .in3(N__11268),
            .lcout(ufifo_utb_txdata_m0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNINUN11_LC_2_9_2 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNINUN11_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNINUN11_LC_2_9_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNINUN11_LC_2_9_2  (
            .in0(N__11269),
            .in1(N__8308),
            .in2(_gnd_net_),
            .in3(N__13377),
            .lcout(ufifo_utb_txdata_m0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNI6GJD2_0_LC_2_9_4 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNI6GJD2_0_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNI6GJD2_0_LC_2_9_4 .LUT_INIT=16'b1011001011110000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNI6GJD2_0_LC_2_9_4  (
            .in0(N__11394),
            .in1(N__9941),
            .in2(N__8302),
            .in3(N__11473),
            .lcout(utb_txdata_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_2_LC_2_9_6 .C_ON=1'b0;
    defparam \resetGen.escKey_2_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_2_LC_2_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.escKey_2_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__11921),
            .in2(_gnd_net_),
            .in3(N__13376),
            .lcout(Lab_UT_dk_de_cr_2_reti),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI9JC39_1_LC_2_9_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI9JC39_1_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI9JC39_1_LC_2_9_7 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI9JC39_1_LC_2_9_7  (
            .in0(N__12179),
            .in1(N__12105),
            .in2(_gnd_net_),
            .in3(N__12040),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_4_LC_2_10_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_2_10_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_2_10_0 .LUT_INIT=16'b1111000010111011;
    LogicCell40 \buart.Z_tx.shifter_4_LC_2_10_0  (
            .in0(N__8272),
            .in1(N__9066),
            .in2(N__8383),
            .in3(N__12042),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22656),
            .ce(N__8372),
            .sr(N__18068));
    defparam \buart.Z_tx.shifter_3_LC_2_10_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_2_10_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_2_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \buart.Z_tx.shifter_3_LC_2_10_1  (
            .in0(N__12041),
            .in1(N__8419),
            .in2(_gnd_net_),
            .in3(N__9019),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22656),
            .ce(N__8372),
            .sr(N__18068));
    defparam \buart.Z_tx.shifter_5_LC_2_10_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_2_10_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_2_10_6 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \buart.Z_tx.shifter_5_LC_2_10_6  (
            .in0(N__8404),
            .in1(N__9067),
            .in2(N__8395),
            .in3(N__12043),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22656),
            .ce(N__8372),
            .sr(N__18068));
    defparam \Lab_UT.scdp.u2.q_esr_1_LC_2_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_1_LC_2_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_1_LC_2_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_1_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15782),
            .lcout(\Lab_UT.scdp.u2.byteToEncrypt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22651),
            .ce(N__8971),
            .sr(N__18039));
    defparam \Lab_UT.scdp.u2.q_esr_2_LC_2_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_2_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_2_LC_2_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_2_LC_2_11_1  (
            .in0(N__15687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scdp.u2.byteToEncrypt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22651),
            .ce(N__8971),
            .sr(N__18039));
    defparam \Lab_UT.scdp.u2.q_esr_3_LC_2_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_3_LC_2_11_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_3_LC_2_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_3_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11934),
            .lcout(\Lab_UT.scdp.byteToEncrypt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22651),
            .ce(N__8971),
            .sr(N__18039));
    defparam \Lab_UT.scdp.u2.q_esr_4_LC_2_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_4_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_4_LC_2_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_4_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13378),
            .lcout(\Lab_UT.scdp.byteToEncrypt_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22651),
            .ce(N__8971),
            .sr(N__18039));
    defparam \Lab_UT.scdp.u2.q_esr_5_LC_2_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_5_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_5_LC_2_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_5_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13438),
            .lcout(\Lab_UT.scdp.u2.byteToEncryptZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22651),
            .ce(N__8971),
            .sr(N__18039));
    defparam \Lab_UT.scdp.u2.q_esr_6_LC_2_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_6_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_6_LC_2_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_6_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17075),
            .lcout(\Lab_UT.scdp.byteToEncrypt_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22651),
            .ce(N__8971),
            .sr(N__18039));
    defparam \Lab_UT.scdp.u2.q_esr_7_LC_2_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_7_LC_2_11_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_7_LC_2_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_7_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16965),
            .lcout(\Lab_UT.scdp.byteToEncrypt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22651),
            .ce(N__8971),
            .sr(N__18039));
    defparam \Lab_UT.scdp.u2.q_esr_0_LC_2_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_0_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_0_LC_2_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_0_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16167),
            .lcout(\Lab_UT.scdp.u2.byteToEncrypt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22651),
            .ce(N__8971),
            .sr(N__18039));
    defparam \Lab_UT.scdp.u2.q_esr_RNIT8JT_0_LC_2_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_RNIT8JT_0_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u2.q_esr_RNIT8JT_0_LC_2_12_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_RNIT8JT_0_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__8446),
            .in2(_gnd_net_),
            .in3(N__9270),
            .lcout(\Lab_UT.scdp.d2eData_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.rdaddr_0_LC_4_1_0 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_0_LC_4_1_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_0_LC_4_1_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_0_LC_4_1_0  (
            .in0(_gnd_net_),
            .in1(N__8516),
            .in2(N__10027),
            .in3(N__10023),
            .lcout(\ufifo.fifo.rdaddrZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_1_0_),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_0 ),
            .clk(N__22698),
            .ce(),
            .sr(N__18050));
    defparam \ufifo.fifo.rdaddr_1_LC_4_1_1 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_1_LC_4_1_1 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_1_LC_4_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_1_LC_4_1_1  (
            .in0(_gnd_net_),
            .in1(N__9530),
            .in2(_gnd_net_),
            .in3(N__8440),
            .lcout(\ufifo.fifo.rdaddrZ0Z_1 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_0 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_1 ),
            .clk(N__22698),
            .ce(),
            .sr(N__18050));
    defparam \ufifo.fifo.rdaddr_2_LC_4_1_2 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_2_LC_4_1_2 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_2_LC_4_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_2_LC_4_1_2  (
            .in0(_gnd_net_),
            .in1(N__9593),
            .in2(_gnd_net_),
            .in3(N__8437),
            .lcout(\ufifo.fifo.rdaddrZ0Z_2 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_1 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_2 ),
            .clk(N__22698),
            .ce(),
            .sr(N__18050));
    defparam \ufifo.fifo.rdaddr_3_LC_4_1_3 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_3_LC_4_1_3 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_3_LC_4_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_3_LC_4_1_3  (
            .in0(_gnd_net_),
            .in1(N__9653),
            .in2(_gnd_net_),
            .in3(N__8434),
            .lcout(\ufifo.fifo.rdaddrZ0Z_3 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_2 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_3 ),
            .clk(N__22698),
            .ce(),
            .sr(N__18050));
    defparam \ufifo.fifo.rdaddr_4_LC_4_1_4 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_4_LC_4_1_4 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_4_LC_4_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_4_LC_4_1_4  (
            .in0(_gnd_net_),
            .in1(N__9770),
            .in2(_gnd_net_),
            .in3(N__8431),
            .lcout(\ufifo.fifo.rdaddrZ0Z_4 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_3 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_4 ),
            .clk(N__22698),
            .ce(),
            .sr(N__18050));
    defparam \ufifo.fifo.rdaddr_5_LC_4_1_5 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_5_LC_4_1_5 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_5_LC_4_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_5_LC_4_1_5  (
            .in0(_gnd_net_),
            .in1(N__9710),
            .in2(_gnd_net_),
            .in3(N__8428),
            .lcout(\ufifo.fifo.rdaddrZ0Z_5 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_4 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_5 ),
            .clk(N__22698),
            .ce(),
            .sr(N__18050));
    defparam \ufifo.fifo.rdaddr_6_LC_4_1_6 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_6_LC_4_1_6 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_6_LC_4_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_6_LC_4_1_6  (
            .in0(_gnd_net_),
            .in1(N__8633),
            .in2(_gnd_net_),
            .in3(N__8425),
            .lcout(\ufifo.fifo.rdaddrZ0Z_6 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_5 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_6 ),
            .clk(N__22698),
            .ce(),
            .sr(N__18050));
    defparam \ufifo.fifo.rdaddr_7_LC_4_1_7 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_7_LC_4_1_7 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_7_LC_4_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_7_LC_4_1_7  (
            .in0(_gnd_net_),
            .in1(N__8693),
            .in2(_gnd_net_),
            .in3(N__8422),
            .lcout(\ufifo.fifo.rdaddrZ0Z_7 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_6 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_7 ),
            .clk(N__22698),
            .ce(),
            .sr(N__18050));
    defparam \ufifo.fifo.rdaddr_8_LC_4_2_0 .C_ON=1'b0;
    defparam \ufifo.fifo.rdaddr_8_LC_4_2_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_8_LC_4_2_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ufifo.fifo.rdaddr_8_LC_4_2_0  (
            .in0(_gnd_net_),
            .in1(N__8579),
            .in2(_gnd_net_),
            .in3(N__8470),
            .lcout(\ufifo.fifo.rdaddrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22694),
            .ce(),
            .sr(N__18047));
    defparam \ufifo.fifo.wraddr_0_LC_4_3_0 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_0_LC_4_3_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_0_LC_4_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_0_LC_4_3_0  (
            .in0(_gnd_net_),
            .in1(N__8606),
            .in2(N__11090),
            .in3(N__11083),
            .lcout(\ufifo.fifo.wraddrZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_3_0_),
            .carryout(\ufifo.fifo.un1_wraddr_cry_0 ),
            .clk(N__22691),
            .ce(),
            .sr(N__18045));
    defparam \ufifo.fifo.wraddr_1_LC_4_3_1 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_1_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_1_LC_4_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_1_LC_4_3_1  (
            .in0(_gnd_net_),
            .in1(N__9567),
            .in2(_gnd_net_),
            .in3(N__8467),
            .lcout(\ufifo.fifo.wraddrZ0Z_1 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_0 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_1 ),
            .clk(N__22691),
            .ce(),
            .sr(N__18045));
    defparam \ufifo.fifo.wraddr_2_LC_4_3_2 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_2_LC_4_3_2 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_2_LC_4_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_2_LC_4_3_2  (
            .in0(_gnd_net_),
            .in1(N__9681),
            .in2(_gnd_net_),
            .in3(N__8464),
            .lcout(\ufifo.fifo.wraddrZ0Z_2 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_1 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_2 ),
            .clk(N__22691),
            .ce(),
            .sr(N__18045));
    defparam \ufifo.fifo.wraddr_3_LC_4_3_3 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_3_LC_4_3_3 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_3_LC_4_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_3_LC_4_3_3  (
            .in0(_gnd_net_),
            .in1(N__9623),
            .in2(_gnd_net_),
            .in3(N__8461),
            .lcout(\ufifo.fifo.wraddrZ0Z_3 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_2 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_3 ),
            .clk(N__22691),
            .ce(),
            .sr(N__18045));
    defparam \ufifo.fifo.wraddr_4_LC_4_3_4 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_4_LC_4_3_4 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_4_LC_4_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_4_LC_4_3_4  (
            .in0(_gnd_net_),
            .in1(N__9798),
            .in2(_gnd_net_),
            .in3(N__8458),
            .lcout(\ufifo.fifo.wraddrZ0Z_4 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_3 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_4 ),
            .clk(N__22691),
            .ce(),
            .sr(N__18045));
    defparam \ufifo.fifo.wraddr_5_LC_4_3_5 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_5_LC_4_3_5 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_5_LC_4_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_5_LC_4_3_5  (
            .in0(_gnd_net_),
            .in1(N__9740),
            .in2(_gnd_net_),
            .in3(N__8455),
            .lcout(\ufifo.fifo.wraddrZ0Z_5 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_4 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_5 ),
            .clk(N__22691),
            .ce(),
            .sr(N__18045));
    defparam \ufifo.fifo.wraddr_6_LC_4_3_6 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_6_LC_4_3_6 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_6_LC_4_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_6_LC_4_3_6  (
            .in0(_gnd_net_),
            .in1(N__8723),
            .in2(_gnd_net_),
            .in3(N__8452),
            .lcout(\ufifo.fifo.wraddrZ0Z_6 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_5 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_6 ),
            .clk(N__22691),
            .ce(),
            .sr(N__18045));
    defparam \ufifo.fifo.wraddr_7_LC_4_3_7 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_7_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_7_LC_4_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_7_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(N__8663),
            .in2(_gnd_net_),
            .in3(N__8449),
            .lcout(\ufifo.fifo.wraddrZ0Z_7 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_6 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_7 ),
            .clk(N__22691),
            .ce(),
            .sr(N__18045));
    defparam \ufifo.fifo.wraddr_8_LC_4_4_0 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_8_LC_4_4_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_8_LC_4_4_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ufifo.fifo.wraddr_8_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__8555),
            .in2(_gnd_net_),
            .in3(N__8740),
            .lcout(\ufifo.fifo.wraddrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22684),
            .ce(),
            .sr(N__18043));
    defparam \resetGen.uu0.counter_gen_label_3__un23_ci_LC_4_5_0 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_3__un23_ci_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_3__un23_ci_LC_4_5_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_3__un23_ci_LC_4_5_0  (
            .in0(N__8480),
            .in1(N__8495),
            .in2(_gnd_net_),
            .in3(N__8816),
            .lcout(\resetGen.un23_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_4_5_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_4_5_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_4_5_1 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \resetGen.reset_count_0_LC_4_5_1  (
            .in0(N__8496),
            .in1(N__22764),
            .in2(_gnd_net_),
            .in3(N__8783),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22677),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_2__un12_ci_LC_4_5_2 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_2__un12_ci_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_2__un12_ci_LC_4_5_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_2__un12_ci_LC_4_5_2  (
            .in0(N__8481),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8494),
            .lcout(\resetGen.un12_ci ),
            .ltout(\resetGen.un12_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_4_5_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_4_5_3 .LUT_INIT=16'b0000000010011010;
    LogicCell40 \resetGen.reset_count_2_LC_4_5_3  (
            .in0(N__8817),
            .in1(N__22763),
            .in2(N__8737),
            .in3(N__8784),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22677),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_RNI8A8U_6_LC_4_5_4 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNI8A8U_6_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNI8A8U_6_LC_4_5_4 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \ufifo.fifo.wraddr_RNI8A8U_6_LC_4_5_4  (
            .in0(N__8727),
            .in1(N__8697),
            .in2(N__8670),
            .in3(N__8634),
            .lcout(\ufifo.fifo.un1_emptyB_NE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_RNIUV7U_8_LC_4_5_5 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNIUV7U_8_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNIUV7U_8_LC_4_5_5 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \ufifo.fifo.wraddr_RNIUV7U_8_LC_4_5_5  (
            .in0(N__8607),
            .in1(N__8580),
            .in2(N__8556),
            .in3(N__8517),
            .lcout(\ufifo.fifo.un1_emptyB_NE_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_10_LC_4_5_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_10_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_10_LC_4_5_6 .LUT_INIT=16'b1100111111011111;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_10_LC_4_5_6  (
            .in0(N__18441),
            .in1(N__18946),
            .in2(N__17615),
            .in3(N__20098),
            .lcout(\Lab_UT.scctrl.g0_7_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_4_5_7 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_4_5_7 .LUT_INIT=16'b0000110000000110;
    LogicCell40 \resetGen.reset_count_1_LC_4_5_7  (
            .in0(N__8497),
            .in1(N__8482),
            .in2(N__8788),
            .in3(N__22765),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22677),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNI56C1D_0_LC_4_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNI56C1D_0_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNI56C1D_0_LC_4_6_1 .LUT_INIT=16'b1111111101100110;
    LogicCell40 \Lab_UT.scdp.u1.q_RNI56C1D_0_LC_4_6_1  (
            .in0(N__9853),
            .in1(N__9271),
            .in2(_gnd_net_),
            .in3(N__9382),
            .lcout(),
            .ltout(\Lab_UT.scdp.q_RNI56C1D_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_0_LC_4_6_2 .C_ON=1'b0;
    defparam \ufifo.txdataD_0_LC_4_6_2 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_0_LC_4_6_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ufifo.txdataD_0_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__8899),
            .in2(N__8836),
            .in3(N__17838),
            .lcout(\ufifo.txdataDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22672),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIQOQA1_0_3_LC_4_6_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_0_3_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_0_3_LC_4_6_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \buart.Z_tx.bitcount_RNIQOQA1_0_3_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(N__11432),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buart__tx_uart_busy_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_6_LC_4_6_4 .C_ON=1'b0;
    defparam \ufifo.txdataD_6_LC_4_6_4 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_6_LC_4_6_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ufifo.txdataD_6_LC_4_6_4  (
            .in0(N__8908),
            .in1(N__17839),
            .in2(_gnd_net_),
            .in3(N__9223),
            .lcout(\ufifo.txdataDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22672),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNO_0_4_LC_4_6_5 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_4_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_4_LC_4_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.reset_count_RNO_0_4_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(N__8748),
            .in2(_gnd_net_),
            .in3(N__8818),
            .lcout(),
            .ltout(\resetGen.reset_count_2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_4_6_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_4_6_6 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_4_6_6 .LUT_INIT=16'b0101010001000100;
    LogicCell40 \resetGen.reset_count_4_LC_4_6_6  (
            .in0(N__8781),
            .in1(N__22744),
            .in2(N__8803),
            .in3(N__8800),
            .lcout(rst_i_3_reti),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22672),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_4_6_7 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_4_6_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_4_6_7 .LUT_INIT=16'b0000000011000110;
    LogicCell40 \resetGen.reset_count_3_LC_4_6_7  (
            .in0(N__8794),
            .in1(N__8749),
            .in2(N__22766),
            .in3(N__8782),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22672),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_3_LC_4_7_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_3_LC_4_7_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.next_state_3_LC_4_7_0 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \Lab_UT.scctrl.next_state_3_LC_4_7_0  (
            .in0(N__21546),
            .in1(N__21489),
            .in2(N__20272),
            .in3(N__14545),
            .lcout(\Lab_UT.scctrl.next_state_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22665),
            .ce(N__14793),
            .sr(N__18071));
    defparam \Lab_UT.scdp.lsBitsi.q_esr_RNI0TMA_3_LC_4_7_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_RNI0TMA_3_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_RNI0TMA_3_LC_4_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_esr_RNI0TMA_3_LC_4_7_1  (
            .in0(N__9148),
            .in1(N__12208),
            .in2(_gnd_net_),
            .in3(N__18164),
            .lcout(\Lab_UT.scdp.lsBitsi.q_esr_RNI0TMAZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNIF1M8_6_LC_4_7_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNIF1M8_6_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNIF1M8_6_LC_4_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNIF1M8_6_LC_4_7_2  (
            .in0(N__18165),
            .in1(N__8881),
            .in2(_gnd_net_),
            .in3(N__9121),
            .lcout(\Lab_UT.scdp.msBitsi.q_esr_RNIF1M8Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNIQQ8E_0_LC_4_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNIQQ8E_0_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNIQQ8E_0_LC_4_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNIQQ8E_0_LC_4_7_3  (
            .in0(N__8959),
            .in1(N__12337),
            .in2(_gnd_net_),
            .in3(N__18166),
            .lcout(\Lab_UT.scdp.msBitsi.q_esr_RNIQQ8EZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_4_LC_4_7_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_4_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_4_LC_4_7_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOP0V3_4_LC_4_7_5  (
            .in0(_gnd_net_),
            .in1(N__10197),
            .in2(_gnd_net_),
            .in3(N__20808),
            .lcout(\buart.Z_rx.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_0_0_LC_4_7_6 .C_ON=1'b0;
    defparam \resetGen.escKey_0_0_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_0_0_LC_4_7_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \resetGen.escKey_0_0_LC_4_7_6  (
            .in0(N__16774),
            .in1(N__15695),
            .in2(_gnd_net_),
            .in3(N__16943),
            .lcout(\resetGen.escKey_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_2_LC_4_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_2_LC_4_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_2_LC_4_8_0 .LUT_INIT=16'b0011001011001000;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_2_LC_4_8_0  (
            .in0(N__8927),
            .in1(N__9109),
            .in2(N__8938),
            .in3(N__8855),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsD_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22657),
            .ce(N__13200),
            .sr(N__18038));
    defparam \Lab_UT.scdp.msBitsi.q_esr_6_LC_4_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_6_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_6_LC_4_8_1 .LUT_INIT=16'b0011001100010010;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_6_LC_4_8_1  (
            .in0(N__9107),
            .in1(N__12259),
            .in2(N__8860),
            .in3(N__8928),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsD_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22657),
            .ce(N__13200),
            .sr(N__18038));
    defparam \Lab_UT.scdp.msBitsi.q_esr_4_LC_4_8_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_4_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_4_LC_4_8_2 .LUT_INIT=16'b1111010011110001;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_4_LC_4_8_2  (
            .in0(N__8929),
            .in1(N__9108),
            .in2(N__12267),
            .in3(N__8859),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsD_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22657),
            .ce(N__13200),
            .sr(N__18038));
    defparam \Lab_UT.scdp.u2.q_esr_RNIKRG71_5_LC_4_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_RNIKRG71_5_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u2.q_esr_RNIKRG71_5_LC_4_8_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_RNIKRG71_5_LC_4_8_3  (
            .in0(N__8875),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10852),
            .lcout(\Lab_UT.scdp.d2eData_5 ),
            .ltout(\Lab_UT.scdp.d2eData_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_o3_3_LC_4_8_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_o3_3_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_o3_3_LC_4_8_4 .LUT_INIT=16'b1111001111111100;
    LogicCell40 \Lab_UT.scdp.b2a0.asciiHex_2_i_o3_3_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(N__9106),
            .in2(N__8863),
            .in3(N__8854),
            .lcout(\Lab_UT.scdp.N_52 ),
            .ltout(\Lab_UT.scdp.N_52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_0_LC_4_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_0_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_0_LC_4_8_5 .LUT_INIT=16'b0110011010010110;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_0_LC_4_8_5  (
            .in0(N__9445),
            .in1(N__8953),
            .in2(N__8962),
            .in3(N__12263),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22657),
            .ce(N__13200),
            .sr(N__18038));
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_0_a2_0_o2_0_LC_4_8_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_0_a2_0_o2_0_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_0_a2_0_o2_0_LC_4_8_6 .LUT_INIT=16'b1101110111101110;
    LogicCell40 \Lab_UT.scdp.b2a0.asciiHex_2_0_a2_0_o2_0_LC_4_8_6  (
            .in0(N__8952),
            .in1(N__12258),
            .in2(_gnd_net_),
            .in3(N__9444),
            .lcout(\Lab_UT.scdp.b2a0.N_55 ),
            .ltout(\Lab_UT.scdp.b2a0.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_1_LC_4_8_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_1_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_1_LC_4_8_7 .LUT_INIT=16'b1100001100000000;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_1_LC_4_8_7  (
            .in0(_gnd_net_),
            .in1(N__8926),
            .in2(N__8914),
            .in3(N__12219),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsD_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22657),
            .ce(N__13200),
            .sr(N__18038));
    defparam \Lab_UT.scctrl.g0_17_N_2L1_LC_4_9_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.g0_17_N_2L1_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.g0_17_N_2L1_LC_4_9_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.scctrl.g0_17_N_2L1_LC_4_9_0  (
            .in0(N__10599),
            .in1(N__12424),
            .in2(N__16505),
            .in3(N__10650),
            .lcout(\Lab_UT.scctrl.g0_17_N_2LZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_fast_RNI1CIH1_2_LC_4_9_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_RNI1CIH1_2_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_0_fast_RNI1CIH1_2_LC_4_9_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \buart.Z_rx.shifter_0_fast_RNI1CIH1_2_LC_4_9_1  (
            .in0(N__12423),
            .in1(N__10649),
            .in2(N__16504),
            .in3(N__10598),
            .lcout(\buart.Z_rx.shifter_0_fast_RNI1CIH1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_fast_2_LC_4_9_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_2_LC_4_9_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_2_LC_4_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_fast_2_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11925),
            .lcout(buart__rx_shifter_0_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22652),
            .ce(N__16752),
            .sr(N__18072));
    defparam \buart.Z_rx.shifter_ret_1_LC_4_9_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_1_LC_4_9_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_1_LC_4_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_1_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15694),
            .lcout(bu_rx_data_i_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22652),
            .ce(N__16752),
            .sr(N__18072));
    defparam \Lab_UT.scdp.a2b.val_0_0_3_LC_4_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_0_0_3_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_0_0_3_LC_4_9_5 .LUT_INIT=16'b0000000101000000;
    LogicCell40 \Lab_UT.scdp.a2b.val_0_0_3_LC_4_9_5  (
            .in0(N__11923),
            .in1(N__16169),
            .in2(N__15704),
            .in3(N__14845),
            .lcout(),
            .ltout(\Lab_UT.scdp.a2b.val_0_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.val_0_3_LC_4_9_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_0_3_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_0_3_LC_4_9_6 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \Lab_UT.scdp.a2b.val_0_3_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__11626),
            .in2(N__8911),
            .in3(N__11924),
            .lcout(\Lab_UT.scdp.val_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.val18_1_i_LC_4_9_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val18_1_i_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val18_1_i_LC_4_9_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \Lab_UT.scdp.a2b.val18_1_i_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(N__16168),
            .in2(_gnd_net_),
            .in3(N__14844),
            .lcout(N_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIM7051_14_LC_4_10_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIM7051_14_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIM7051_14_LC_4_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIM7051_14_LC_4_10_0  (
            .in0(N__10840),
            .in1(N__10677),
            .in2(N__11797),
            .in3(N__11824),
            .lcout(\Lab_UT.scdp.d2eData_3_6 ),
            .ltout(\Lab_UT.scdp.d2eData_3_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_esr_RNIA29D1_2_LC_4_10_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_esr_RNIA29D1_2_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_esr_RNIA29D1_2_LC_4_10_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \Lab_UT.scdp.u0.q_esr_RNIA29D1_2_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9091),
            .in3(N__9088),
            .lcout(\Lab_UT.scdp.e2dData_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_esr_2_LC_4_10_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_esr_2_LC_4_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u0.q_esr_2_LC_4_10_2 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \Lab_UT.scdp.u0.q_esr_2_LC_4_10_2  (
            .in0(N__15696),
            .in1(N__15772),
            .in2(_gnd_net_),
            .in3(N__15818),
            .lcout(\Lab_UT.scdp.u0.byteToDecrypt_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22645),
            .ce(N__13126),
            .sr(N__18040));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2_0_LC_4_10_4 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2_0_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2_0_LC_4_10_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2_0_LC_4_10_4  (
            .in0(N__11395),
            .in1(N__9942),
            .in2(_gnd_net_),
            .in3(N__11468),
            .lcout(),
            .ltout(\ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIR7FP3_0_LC_4_10_5 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIR7FP3_0_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIR7FP3_0_LC_4_10_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIR7FP3_0_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(N__9082),
            .in2(N__9070),
            .in3(N__9065),
            .lcout(utb_txdata_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_1_LC_4_11_0 .C_ON=1'b0;
    defparam \ufifo.txdataD_1_LC_4_11_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_1_LC_4_11_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ufifo.txdataD_1_LC_4_11_0  (
            .in0(N__8989),
            .in1(N__17830),
            .in2(_gnd_net_),
            .in3(N__9178),
            .lcout(\ufifo.txdataDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22639),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8_1_LC_4_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8_1_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8_1_LC_4_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8_1_LC_4_11_1  (
            .in0(N__8998),
            .in1(N__9154),
            .in2(_gnd_net_),
            .in3(N__18155),
            .lcout(\Lab_UT.scdp.msBitsi.q_esr_RNI5NL8Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_5_LC_4_11_2 .C_ON=1'b0;
    defparam \ufifo.txdataD_5_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_5_LC_4_11_2 .LUT_INIT=16'b1111001111100010;
    LogicCell40 \ufifo.txdataD_5_LC_4_11_2  (
            .in0(N__9381),
            .in1(N__17832),
            .in2(N__13156),
            .in3(N__11191),
            .lcout(\ufifo.txdataDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22639),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u2.q_esr_ctle_7_LC_4_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_ctle_7_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u2.q_esr_ctle_7_LC_4_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_ctle_7_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(N__18091),
            .in2(_gnd_net_),
            .in3(N__12823),
            .lcout(\Lab_UT.scdp.u2.sccEldByte_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI7PL8_2_LC_4_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI7PL8_2_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI7PL8_2_LC_4_11_4 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNI7PL8_2_LC_4_11_4  (
            .in0(N__18156),
            .in1(_gnd_net_),
            .in2(N__9301),
            .in3(N__9208),
            .lcout(),
            .ltout(\Lab_UT.scdp.msBitsi.L4_tx_data_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_2_LC_4_11_5 .C_ON=1'b0;
    defparam \ufifo.txdataD_2_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_2_LC_4_11_5 .LUT_INIT=16'b0000101001001110;
    LogicCell40 \ufifo.txdataD_2_LC_4_11_5  (
            .in0(N__17831),
            .in1(N__9487),
            .in2(N__9196),
            .in3(N__9380),
            .lcout(\ufifo.txdataDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22639),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNID22R_1_LC_4_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNID22R_1_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNID22R_1_LC_4_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNID22R_1_LC_4_11_6  (
            .in0(N__10737),
            .in1(N__10689),
            .in2(N__10813),
            .in3(N__12526),
            .lcout(\Lab_UT.scdp.d2eData_3_1 ),
            .ltout(\Lab_UT.scdp.d2eData_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNIABC1D_1_LC_4_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNIABC1D_1_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNIABC1D_1_LC_4_11_7 .LUT_INIT=16'b1111111100111100;
    LogicCell40 \Lab_UT.scdp.u1.q_RNIABC1D_1_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(N__14002),
            .in2(N__9181),
            .in3(N__9379),
            .lcout(\Lab_UT.scdp.q_RNIABC1D_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u2.q_esr_RNI2EJT_1_LC_4_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_RNI2EJT_1_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u2.q_esr_RNI2EJT_1_LC_4_12_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_RNI2EJT_1_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(N__9172),
            .in2(_gnd_net_),
            .in3(N__9291),
            .lcout(\Lab_UT.scdp.d2eData_1 ),
            .ltout(\Lab_UT.scdp.d2eData_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.b2a1.lowerTen_LC_4_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a1.lowerTen_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a1.lowerTen_LC_4_12_1 .LUT_INIT=16'b0110011001100000;
    LogicCell40 \Lab_UT.scdp.b2a1.lowerTen_LC_4_12_1  (
            .in0(N__9137),
            .in1(N__9401),
            .in2(N__9160),
            .in3(N__9326),
            .lcout(\Lab_UT.scdp.lsBits_6 ),
            .ltout(\Lab_UT.scdp.lsBits_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lsBitsi.q_esr_1_LC_4_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_1_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_1_LC_4_12_2 .LUT_INIT=16'b1100110000111100;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_esr_1_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(N__9311),
            .in2(N__9157),
            .in3(N__12356),
            .lcout(\Lab_UT.scdp.lsBitsD_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22633),
            .ce(N__13204),
            .sr(N__18042));
    defparam \Lab_UT.scdp.lsBitsi.q_esr_3_LC_4_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_3_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_3_LC_4_12_3 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_esr_3_LC_4_12_3  (
            .in0(N__9138),
            .in1(N__9402),
            .in2(_gnd_net_),
            .in3(N__12304),
            .lcout(\Lab_UT.scdp.lsBitsi.lsBitsD_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22633),
            .ce(N__13204),
            .sr(N__18042));
    defparam \Lab_UT.scdp.lsBitsi.q_esr_6_LC_4_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_6_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_6_LC_4_12_4 .LUT_INIT=16'b0110011001100000;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_esr_6_LC_4_12_4  (
            .in0(N__9403),
            .in1(N__9139),
            .in2(N__9331),
            .in3(N__9315),
            .lcout(\Lab_UT.scdp.lsBitsD_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22633),
            .ce(N__13204),
            .sr(N__18042));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIO7U41_10_LC_4_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIO7U41_10_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIO7U41_10_LC_4_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIO7U41_10_LC_4_12_5  (
            .in0(N__10824),
            .in1(N__10725),
            .in2(N__10915),
            .in3(N__11779),
            .lcout(\Lab_UT.scdp.d2eData_3_2 ),
            .ltout(\Lab_UT.scdp.d2eData_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u2.q_esr_RNIEKF71_2_LC_4_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_RNIEKF71_2_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u2.q_esr_RNIEKF71_2_LC_4_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_RNIEKF71_2_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9346),
            .in3(N__9343),
            .lcout(\Lab_UT.scdp.d2eData_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lsBitsi.q_esr_2_LC_4_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_2_LC_4_12_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_2_LC_4_12_7 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_esr_2_LC_4_12_7  (
            .in0(N__12357),
            .in1(N__9327),
            .in2(N__9316),
            .in3(N__12305),
            .lcout(\Lab_UT.scdp.lsBitsD_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22633),
            .ce(N__13204),
            .sr(N__18042));
    defparam \Lab_UT.scdp.pinst0.un12_pValid_0_LC_4_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.pinst0.un12_pValid_0_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.pinst0.un12_pValid_0_LC_4_13_0 .LUT_INIT=16'b0001010000101000;
    LogicCell40 \Lab_UT.scdp.pinst0.un12_pValid_0_LC_4_13_0  (
            .in0(N__9849),
            .in1(N__9292),
            .in2(N__14001),
            .in3(N__9257),
            .lcout(),
            .ltout(\Lab_UT.scdp.pinst0.un12_pValidZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.pinst0.un12_pValid_LC_4_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.pinst0.un12_pValid_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.pinst0.un12_pValid_LC_4_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scdp.pinst0.un12_pValid_LC_4_13_1  (
            .in0(N__9460),
            .in1(N__11183),
            .in2(N__9277),
            .in3(N__9483),
            .lcout(\Lab_UT.scdp.un12_pValid ),
            .ltout(\Lab_UT.scdp.un12_pValid_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.pinst0.pValid_LC_4_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.pinst0.pValid_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.pinst0.pValid_LC_4_13_2 .LUT_INIT=16'b1111001101110111;
    LogicCell40 \Lab_UT.scdp.pinst0.pValid_LC_4_13_2  (
            .in0(N__11184),
            .in1(N__9471),
            .in2(N__9274),
            .in3(N__9234),
            .lcout(\Lab_UT.scdp.pValid_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI9U1R_0_LC_4_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI9U1R_0_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI9U1R_0_LC_4_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI9U1R_0_LC_4_13_3  (
            .in0(N__10768),
            .in1(N__10926),
            .in2(N__11013),
            .in3(N__12544),
            .lcout(\Lab_UT.scdp.d2eData_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNIDHFGA_3_LC_4_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNIDHFGA_3_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNIDHFGA_3_LC_4_13_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.scdp.u0.q_RNIDHFGA_3_LC_4_13_4  (
            .in0(N__9472),
            .in1(N__9241),
            .in2(_gnd_net_),
            .in3(N__9235),
            .lcout(\Lab_UT.scdp.q_RNIDHFGA_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_esr_RNIDBBI1_2_LC_4_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_esr_RNIDBBI1_2_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_esr_RNIDBBI1_2_LC_4_13_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.scdp.u1.q_esr_RNIDBBI1_2_LC_4_13_5  (
            .in0(N__9214),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12625),
            .lcout(\Lab_UT.scdp.e2dData_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNITJGS_3_LC_4_13_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNITJGS_3_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNITJGS_3_LC_4_13_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.u0.q_RNITJGS_3_LC_4_13_7  (
            .in0(N__10949),
            .in1(N__11040),
            .in2(N__10797),
            .in3(N__11160),
            .lcout(\Lab_UT.scdp.N_59_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.pinst0.un12_pValid_1_LC_4_14_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.pinst0.un12_pValid_1_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.pinst0.un12_pValid_1_LC_4_14_0 .LUT_INIT=16'b0001010000101000;
    LogicCell40 \Lab_UT.scdp.pinst0.un12_pValid_1_LC_4_14_0  (
            .in0(N__9824),
            .in1(N__9438),
            .in2(N__11848),
            .in3(N__9393),
            .lcout(\Lab_UT.scdp.pinst0.un12_pValidZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI239E_4_LC_4_14_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI239E_4_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI239E_4_LC_4_14_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNI239E_4_LC_4_14_1  (
            .in0(N__12286),
            .in1(N__9454),
            .in2(_gnd_net_),
            .in3(N__18141),
            .lcout(\Lab_UT.scdp.msBitsi.q_esr_RNI239EZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIN7V41_4_LC_4_14_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIN7V41_4_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIN7V41_4_LC_4_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIN7V41_4_LC_4_14_2  (
            .in0(N__11758),
            .in1(N__10980),
            .in2(N__10969),
            .in3(N__12508),
            .lcout(\Lab_UT.scdp.d2eData_3_4 ),
            .ltout(\Lab_UT.scdp.d2eData_3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNIIAV0D_0_LC_4_14_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNIIAV0D_0_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNIIAV0D_0_LC_4_14_3 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \Lab_UT.scdp.u0.q_RNIIAV0D_0_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__11847),
            .in2(N__9427),
            .in3(N__9374),
            .lcout(),
            .ltout(\Lab_UT.scdp.q_RNIIAV0D_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_4_LC_4_14_4 .C_ON=1'b0;
    defparam \ufifo.txdataD_4_LC_4_14_4 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_4_LC_4_14_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ufifo.txdataD_4_LC_4_14_4  (
            .in0(N__17842),
            .in1(_gnd_net_),
            .in2(N__9424),
            .in3(N__9421),
            .lcout(\ufifo.txdataDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22625),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNISBU41_3_LC_4_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNISBU41_3_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNISBU41_3_LC_4_14_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNISBU41_3_LC_4_14_5  (
            .in0(N__10753),
            .in1(N__11724),
            .in2(N__10900),
            .in3(N__10996),
            .lcout(\Lab_UT.scdp.d2eData_3_3 ),
            .ltout(\Lab_UT.scdp.d2eData_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNIRM8BD_3_LC_4_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNIRM8BD_3_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNIRM8BD_3_LC_4_14_6 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNIRM8BD_3_LC_4_14_6  (
            .in0(N__9375),
            .in1(_gnd_net_),
            .in2(N__9349),
            .in3(N__9825),
            .lcout(),
            .ltout(\Lab_UT.scdp.q_RNIRM8BD_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_3_LC_4_14_7 .C_ON=1'b0;
    defparam \ufifo.txdataD_3_LC_4_14_7 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_3_LC_4_14_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ufifo.txdataD_3_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(N__9880),
            .in2(N__9871),
            .in3(N__17841),
            .lcout(\ufifo.txdataDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22625),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_0_LC_4_15_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_0_LC_4_15_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u1.q_0_LC_4_15_0 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \Lab_UT.scdp.u1.q_0_LC_4_15_0  (
            .in0(N__11869),
            .in1(N__14019),
            .in2(_gnd_net_),
            .in3(N__9848),
            .lcout(\Lab_UT.scdp.byteToDecrypt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22620),
            .ce(),
            .sr(N__18049));
    defparam \Lab_UT.scdp.u1.q_3_LC_4_15_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_3_LC_4_15_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u1.q_3_LC_4_15_5 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \Lab_UT.scdp.u1.q_3_LC_4_15_5  (
            .in0(N__14020),
            .in1(N__11148),
            .in2(_gnd_net_),
            .in3(N__9826),
            .lcout(\Lab_UT.scdp.byteToDecrypt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22620),
            .ce(),
            .sr(N__18049));
    defparam \ufifo.fifo.wraddr_RNI028U_4_LC_5_3_0 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNI028U_4_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNI028U_4_LC_5_3_0 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \ufifo.fifo.wraddr_RNI028U_4_LC_5_3_0  (
            .in0(N__9797),
            .in1(N__9774),
            .in2(N__9744),
            .in3(N__9714),
            .lcout(\ufifo.fifo.un1_emptyB_NE_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_RNIOP7U_2_LC_5_3_2 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNIOP7U_2_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNIOP7U_2_LC_5_3_2 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \ufifo.fifo.wraddr_RNIOP7U_2_LC_5_3_2  (
            .in0(N__9680),
            .in1(N__9657),
            .in2(N__9627),
            .in3(N__9597),
            .lcout(),
            .ltout(\ufifo.fifo.un1_emptyB_NE_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_RNIHJBD1_1_LC_5_3_3 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNIHJBD1_1_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNIHJBD1_1_LC_5_3_3 .LUT_INIT=16'b1100000000110000;
    LogicCell40 \ufifo.fifo.wraddr_RNIHJBD1_1_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__9566),
            .in2(N__9547),
            .in3(N__9537),
            .lcout(\ufifo.fifo.un1_emptyB_NE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIN78A_0_LC_5_3_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIN78A_0_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIN78A_0_LC_5_3_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIN78A_0_LC_5_3_5  (
            .in0(N__18442),
            .in1(N__18953),
            .in2(_gnd_net_),
            .in3(N__20096),
            .lcout(\Lab_UT.scctrl.g0_16_mb_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_5_LC_5_4_0 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_5_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_5_LC_5_4_0 .LUT_INIT=16'b1011101110110000;
    LogicCell40 \ufifo.tx_fsm.cstate_5_LC_5_4_0  (
            .in0(N__11519),
            .in1(N__11301),
            .in2(N__11319),
            .in3(N__11485),
            .lcout(\ufifo.tx_fsm.cstateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22678),
            .ce(),
            .sr(N__9966));
    defparam \ufifo.tx_fsm.cstate_4_LC_5_4_6 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_4_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_4_LC_5_4_6 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \ufifo.tx_fsm.cstate_4_LC_5_4_6  (
            .in0(N__9511),
            .in1(N__11518),
            .in2(_gnd_net_),
            .in3(N__12175),
            .lcout(\ufifo.tx_fsm.cstateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22678),
            .ce(),
            .sr(N__9966));
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_5_5_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_5_5_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_tx.bitcount_RNIQOQA1_3_LC_5_5_0  (
            .in0(N__10134),
            .in1(N__10116),
            .in2(N__10099),
            .in3(N__11964),
            .lcout(buart__tx_uart_busy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_1_LC_5_5_1 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_1_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_1_LC_5_5_1 .LUT_INIT=16'b1010100011111000;
    LogicCell40 \ufifo.tx_fsm.cstate_1_LC_5_5_1  (
            .in0(N__11241),
            .in1(N__16069),
            .in2(N__10042),
            .in3(N__11293),
            .lcout(\ufifo.tx_fsm.cstateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22673),
            .ce(),
            .sr(N__9973));
    defparam \ufifo.fifo.wraddr_RNINV384_1_LC_5_5_2 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNINV384_1_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNINV384_1_LC_5_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ufifo.fifo.wraddr_RNINV384_1_LC_5_5_2  (
            .in0(N__10081),
            .in1(N__10075),
            .in2(N__10066),
            .in3(N__10054),
            .lcout(\ufifo.emptyB_0 ),
            .ltout(\ufifo.emptyB_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNO_0_2_LC_5_5_3 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNO_0_2_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNO_0_2_LC_5_5_3 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \ufifo.tx_fsm.cstate_RNO_0_2_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(N__11517),
            .in2(N__10045),
            .in3(N__11452),
            .lcout(),
            .ltout(\ufifo.tx_fsm.N_62_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_2_LC_5_5_4 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_2_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_2_LC_5_5_4 .LUT_INIT=16'b1111110010101000;
    LogicCell40 \ufifo.tx_fsm.cstate_2_LC_5_5_4  (
            .in0(N__11294),
            .in1(N__10038),
            .in2(N__10030),
            .in3(N__11524),
            .lcout(\ufifo.popFifo ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22673),
            .ce(),
            .sr(N__9973));
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_1_1_LC_5_6_0 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_1_1_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_1_1_LC_5_6_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNO_1_1_LC_5_6_0  (
            .in0(N__9943),
            .in1(N__11370),
            .in2(_gnd_net_),
            .in3(N__20283),
            .lcout(\ufifo.emitcrlf_fsm.cstate_srsts_sn_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_7_0_LC_5_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_7_0_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_7_0_LC_5_6_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_7_0_LC_5_6_1  (
            .in0(N__16163),
            .in1(N__17073),
            .in2(N__15703),
            .in3(N__16960),
            .lcout(\Lab_UT.scctrl.m24_e_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_2_LC_5_6_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_2_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_2_LC_5_6_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIPVCP_2_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__12435),
            .in2(_gnd_net_),
            .in3(N__10657),
            .lcout(),
            .ltout(\buart.Z_rx.bitcountlde_i_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_5_6_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_5_6_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_5_6_3  (
            .in0(N__10490),
            .in1(N__10552),
            .in2(N__9883),
            .in3(N__10608),
            .lcout(\buart.Z_rx.N_58 ),
            .ltout(\buart.Z_rx.N_58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_6_4 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_6_4 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \buart.Z_rx.hh_RNIJ3K62_0_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(N__10714),
            .in2(N__10222),
            .in3(N__10219),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(\buart.Z_rx.startbit_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIELQA6_4_LC_5_6_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIELQA6_4_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIELQA6_4_LC_5_6_5 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIELQA6_4_LC_5_6_5  (
            .in0(N__20787),
            .in1(N__10198),
            .in2(N__10186),
            .in3(N__10183),
            .lcout(\buart.Z_rx.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.g0_17_N_3L3_LC_5_6_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.g0_17_N_3L3_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.g0_17_N_3L3_LC_5_6_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.scctrl.g0_17_N_3L3_LC_5_6_7  (
            .in0(N__14855),
            .in1(N__10486),
            .in2(_gnd_net_),
            .in3(N__10551),
            .lcout(\Lab_UT.scctrl.g0_17_N_3LZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_5_7_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_5_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(N__10603),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_5_7_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_5_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(N__10546),
            .in2(_gnd_net_),
            .in3(N__10147),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_5_7_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_5_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(N__12430),
            .in2(_gnd_net_),
            .in3(N__10144),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_5_7_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_5_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(N__10656),
            .in2(_gnd_net_),
            .in3(N__10141),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_4_LC_5_7_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_4_LC_5_7_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_4_LC_5_7_4 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_4_LC_5_7_4  (
            .in0(N__10357),
            .in1(N__10305),
            .in2(N__10498),
            .in3(N__10138),
            .lcout(buart__rx_bitcount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22658),
            .ce(N__10279),
            .sr(N__18074));
    defparam \buart.Z_rx.bitcount_es_RNIGTPI1_3_LC_5_8_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIGTPI1_3_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIGTPI1_3_LC_5_8_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIGTPI1_3_LC_5_8_0  (
            .in0(N__10647),
            .in1(N__10589),
            .in2(N__10548),
            .in3(N__10477),
            .lcout(\buart.Z_rx.bitcount_es_RNIGTPI1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNI4E361_2_LC_5_8_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNI4E361_2_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNI4E361_2_LC_5_8_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \buart.Z_rx.bitcount_es_RNI4E361_2_LC_5_8_3  (
            .in0(N__10651),
            .in1(N__10534),
            .in2(_gnd_net_),
            .in3(N__12425),
            .lcout(\buart.Z_rx.N_41_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_3_LC_5_8_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_3_LC_5_8_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_3_LC_5_8_4 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_3_LC_5_8_4  (
            .in0(N__10309),
            .in1(N__10360),
            .in2(N__10393),
            .in3(N__10652),
            .lcout(buart__rx_bitcount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22653),
            .ce(N__10278),
            .sr(N__18069));
    defparam \buart.Z_rx.bitcount_es_1_LC_5_8_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_1_LC_5_8_5 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_1_LC_5_8_5 .LUT_INIT=16'b0000111101100110;
    LogicCell40 \buart.Z_rx.bitcount_es_1_LC_5_8_5  (
            .in0(N__10547),
            .in1(N__10384),
            .in2(N__10373),
            .in3(N__10307),
            .lcout(buart__rx_bitcount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22653),
            .ce(N__10278),
            .sr(N__18069));
    defparam \buart.Z_rx.bitcount_es_0_LC_5_8_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_0_LC_5_8_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_0_LC_5_8_6 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_0_LC_5_8_6  (
            .in0(N__10306),
            .in1(N__10359),
            .in2(N__13965),
            .in3(N__10590),
            .lcout(buart__rx_bitcount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22653),
            .ce(N__10278),
            .sr(N__18069));
    defparam \buart.Z_rx.bitcount_es_2_LC_5_8_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_2_LC_5_8_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_2_LC_5_8_7 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_2_LC_5_8_7  (
            .in0(N__10358),
            .in1(N__10308),
            .in2(N__10288),
            .in3(N__12426),
            .lcout(buart__rx_bitcount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22653),
            .ce(N__10278),
            .sr(N__18069));
    defparam \Lab_UT.dk.de_bigL_LC_5_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigL_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigL_LC_5_9_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dk.de_bigL_LC_5_9_0  (
            .in0(N__10249),
            .in1(N__10665),
            .in2(N__10258),
            .in3(N__10420),
            .lcout(\Lab_UT.de_bigL ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.de_bigL_sx_LC_5_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigL_sx_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigL_sx_LC_5_9_1 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \Lab_UT.dk.de_bigL_sx_LC_5_9_1  (
            .in0(N__10494),
            .in1(N__10535),
            .in2(N__14854),
            .in3(N__10591),
            .lcout(\Lab_UT.dk.de_bigL_sxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.de_bigL_3_LC_5_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigL_3_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigL_3_LC_5_9_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dk.de_bigL_3_LC_5_9_2  (
            .in0(N__16549),
            .in1(N__16846),
            .in2(N__11674),
            .in3(N__13474),
            .lcout(\Lab_UT.de_bigL_3 ),
            .ltout(\Lab_UT.de_bigL_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.g0_17_N_4L5_LC_5_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.g0_17_N_4L5_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.g0_17_N_4L5_LC_5_9_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.scctrl.g0_17_N_4L5_LC_5_9_3  (
            .in0(N__10666),
            .in1(N__10243),
            .in2(N__10234),
            .in3(N__10231),
            .lcout(\Lab_UT.scctrl.g0_17_N_4LZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.de_bigL_0_LC_5_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigL_0_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigL_0_LC_5_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dk.de_bigL_0_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(N__17021),
            .in2(_gnd_net_),
            .in3(N__13250),
            .lcout(\Lab_UT.de_bigL_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_ret_3_LC_5_9_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_3_LC_5_9_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_3_LC_5_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_3_LC_5_9_6  (
            .in0(N__17022),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22646),
            .ce(N__16753),
            .sr(N__18075));
    defparam \Lab_UT.dk.de_bigD_1_0_LC_5_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigD_1_0_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigD_1_0_LC_5_9_7 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \Lab_UT.dk.de_bigD_1_0_LC_5_9_7  (
            .in0(N__16489),
            .in1(_gnd_net_),
            .in2(N__12434),
            .in3(N__10648),
            .lcout(\Lab_UT.dk.de_bigD_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_6_LC_5_10_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_6_LC_5_10_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_6_LC_5_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_6_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16854),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22640),
            .ce(N__16754),
            .sr(N__18076));
    defparam \Lab_UT.dk.de_bigD_sx_LC_5_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigD_sx_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigD_sx_LC_5_10_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \Lab_UT.dk.de_bigD_sx_LC_5_10_1  (
            .in0(N__10495),
            .in1(N__10549),
            .in2(N__16899),
            .in3(N__10604),
            .lcout(\Lab_UT.dk.de_bigD_sxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIF6D61_4_LC_5_10_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIF6D61_4_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIF6D61_4_LC_5_10_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIF6D61_4_LC_5_10_2  (
            .in0(N__10550),
            .in1(N__16853),
            .in2(_gnd_net_),
            .in3(N__10496),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_es_RNIF6D61Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_fast_RNI639J4_2_LC_5_10_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_RNI639J4_2_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_0_fast_RNI639J4_2_LC_5_10_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \buart.Z_rx.shifter_0_fast_RNI639J4_2_LC_5_10_3  (
            .in0(N__10444),
            .in1(N__10435),
            .in2(N__10438),
            .in3(N__16433),
            .lcout(shifter_0_fast_RNI639J4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.de_bigD_0_LC_5_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigD_0_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigD_0_LC_5_10_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dk.de_bigD_0_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__16550),
            .in2(_gnd_net_),
            .in3(N__17019),
            .lcout(Lab_UT_dk_de_bigD_0),
            .ltout(Lab_UT_dk_de_bigD_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.de_bigD_LC_5_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigD_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigD_LC_5_10_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dk.de_bigD_LC_5_10_5  (
            .in0(N__10429),
            .in1(N__16432),
            .in2(N__10423),
            .in3(N__10419),
            .lcout(\Lab_UT.de_bigD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_7_LC_5_10_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_7_LC_5_10_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_7_LC_5_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_7_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10710),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22640),
            .ce(N__16754),
            .sr(N__18076));
    defparam \Lab_UT.dk.de_bigE_1_LC_5_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigE_1_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigE_1_LC_5_10_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \Lab_UT.dk.de_bigE_1_LC_5_10_7  (
            .in0(N__17020),
            .in1(_gnd_net_),
            .in2(N__16900),
            .in3(N__16490),
            .lcout(\Lab_UT.dk.de_bigEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_18_LC_5_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_18_LC_5_11_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_18_LC_5_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_18_LC_5_11_0  (
            .in0(N__12738),
            .in1(N__14893),
            .in2(_gnd_net_),
            .in3(N__10690),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22634),
            .ce(N__12469),
            .sr(N__18078));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_23_LC_5_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_23_LC_5_11_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_23_LC_5_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_23_LC_5_11_1  (
            .in0(N__13747),
            .in1(N__10839),
            .in2(_gnd_net_),
            .in3(N__12741),
            .lcout(\Lab_UT.scdp.prng_lfsr_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22634),
            .ce(N__12469),
            .sr(N__18078));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_17_LC_5_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_17_LC_5_11_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_17_LC_5_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_17_LC_5_11_2  (
            .in0(N__12737),
            .in1(N__14929),
            .in2(_gnd_net_),
            .in3(N__10767),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22634),
            .ce(N__12469),
            .sr(N__18078));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_25_LC_5_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_25_LC_5_11_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_25_LC_5_11_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_25_LC_5_11_3  (
            .in0(N__12907),
            .in1(N__11014),
            .in2(_gnd_net_),
            .in3(N__12742),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22634),
            .ce(N__12469),
            .sr(N__18078));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_7_LC_5_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_7_LC_5_11_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_7_LC_5_11_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_7_LC_5_11_4  (
            .in0(N__12739),
            .in1(N__15412),
            .in2(_gnd_net_),
            .in3(N__11819),
            .lcout(\Lab_UT.scdp.prng_lfsr_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22634),
            .ce(N__12469),
            .sr(N__18078));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_14_LC_5_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_14_LC_5_11_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_14_LC_5_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_14_LC_5_11_5  (
            .in0(N__13609),
            .in1(N__12483),
            .in2(_gnd_net_),
            .in3(N__12740),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22634),
            .ce(N__12469),
            .sr(N__18078));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_15_LC_5_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_15_LC_5_11_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_15_LC_5_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_15_LC_5_11_6  (
            .in0(N__12736),
            .in1(N__11125),
            .in2(_gnd_net_),
            .in3(N__10678),
            .lcout(\Lab_UT.scdp.prng_lfsr_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22634),
            .ce(N__12469),
            .sr(N__18078));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_30_LC_5_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_30_LC_5_11_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_30_LC_5_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_30_LC_5_11_7  (
            .in0(N__13816),
            .in1(N__10870),
            .in2(_gnd_net_),
            .in3(N__12743),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22634),
            .ce(N__12469),
            .sr(N__18078));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_22_LC_5_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_22_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_22_LC_5_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_22_LC_5_12_0  (
            .in0(N__12796),
            .in1(N__13855),
            .in2(_gnd_net_),
            .in3(N__10884),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22629),
            .ce(N__12468),
            .sr(N__18080));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_19_LC_5_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_19_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_19_LC_5_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_19_LC_5_12_1  (
            .in0(N__13873),
            .in1(N__10825),
            .in2(_gnd_net_),
            .in3(N__12800),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22629),
            .ce(N__12468),
            .sr(N__18080));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_10_LC_5_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_10_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_10_LC_5_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_10_LC_5_12_2  (
            .in0(N__12795),
            .in1(N__14173),
            .in2(_gnd_net_),
            .in3(N__10738),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22629),
            .ce(N__12468),
            .sr(N__18080));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_4_LC_5_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_4_LC_5_12_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_4_LC_5_12_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_4_LC_5_12_3  (
            .in0(N__15454),
            .in1(N__10752),
            .in2(_gnd_net_),
            .in3(N__12801),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22629),
            .ce(N__12468),
            .sr(N__18080));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_26_LC_5_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_26_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_26_LC_5_12_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_26_LC_5_12_4  (
            .in0(N__12797),
            .in1(_gnd_net_),
            .in2(N__13795),
            .in3(N__10812),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22629),
            .ce(N__12468),
            .sr(N__18080));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_16_LC_5_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_16_LC_5_12_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_16_LC_5_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_16_LC_5_12_5  (
            .in0(N__10790),
            .in1(N__14947),
            .in2(_gnd_net_),
            .in3(N__12799),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22629),
            .ce(N__12468),
            .sr(N__18080));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_3_LC_5_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_3_LC_5_12_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_3_LC_5_12_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_3_LC_5_12_6  (
            .in0(N__12798),
            .in1(N__15052),
            .in2(_gnd_net_),
            .in3(N__11778),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22629),
            .ce(N__12468),
            .sr(N__18080));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_9_LC_5_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_9_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_9_LC_5_12_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_9_LC_5_12_7  (
            .in0(N__12598),
            .in1(N__10927),
            .in2(_gnd_net_),
            .in3(N__12802),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22629),
            .ce(N__12468),
            .sr(N__18080));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_11_LC_5_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_11_LC_5_13_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_11_LC_5_13_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_11_LC_5_13_0  (
            .in0(N__12787),
            .in1(N__11107),
            .in2(_gnd_net_),
            .in3(N__10726),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22626),
            .ce(N__12466),
            .sr(N__18082));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_24_LC_5_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_24_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_24_LC_5_13_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_24_LC_5_13_1  (
            .in0(N__11039),
            .in1(N__12450),
            .in2(_gnd_net_),
            .in3(N__12791),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22626),
            .ce(N__12466),
            .sr(N__18082));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_20_LC_5_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_20_LC_5_13_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_20_LC_5_13_2 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_20_LC_5_13_2  (
            .in0(N__12788),
            .in1(N__10995),
            .in2(N__12864),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22626),
            .ce(N__12466),
            .sr(N__18082));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_28_LC_5_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_28_LC_5_13_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_28_LC_5_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_28_LC_5_13_3  (
            .in0(N__12841),
            .in1(N__10899),
            .in2(_gnd_net_),
            .in3(N__12793),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22626),
            .ce(N__12466),
            .sr(N__18082));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_21_LC_5_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_21_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_21_LC_5_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_21_LC_5_13_4  (
            .in0(N__12789),
            .in1(N__12577),
            .in2(_gnd_net_),
            .in3(N__10981),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22626),
            .ce(N__12466),
            .sr(N__18082));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_29_LC_5_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_29_LC_5_13_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_29_LC_5_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_29_LC_5_13_5  (
            .in0(N__12559),
            .in1(N__10968),
            .in2(_gnd_net_),
            .in3(N__12794),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22626),
            .ce(N__12466),
            .sr(N__18082));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_8_LC_5_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_8_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_8_LC_5_13_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_8_LC_5_13_6  (
            .in0(N__12790),
            .in1(_gnd_net_),
            .in2(N__12886),
            .in3(N__10950),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22626),
            .ce(N__12466),
            .sr(N__18082));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_27_LC_5_13_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_27_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_27_LC_5_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_27_LC_5_13_7  (
            .in0(N__13699),
            .in1(N__10914),
            .in2(_gnd_net_),
            .in3(N__12792),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22626),
            .ce(N__12466),
            .sr(N__18082));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIRBV41_13_LC_5_14_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIRBV41_13_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIRBV41_13_LC_5_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIRBV41_13_LC_5_14_0  (
            .in0(N__10885),
            .in1(N__12484),
            .in2(N__10869),
            .in3(N__11743),
            .lcout(\Lab_UT.scdp.d2eData_3_5 ),
            .ltout(\Lab_UT.scdp.d2eData_3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNI5V781_1_LC_5_14_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNI5V781_1_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNI5V781_1_LC_5_14_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \Lab_UT.scdp.u0.q_RNI5V781_1_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11194),
            .in3(N__11169),
            .lcout(\Lab_UT.scdp.e2dData_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_1_LC_5_14_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_1_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u0.q_1_LC_5_14_2 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \Lab_UT.scdp.u0.q_1_LC_5_14_2  (
            .in0(N__11170),
            .in1(N__14040),
            .in2(_gnd_net_),
            .in3(N__12951),
            .lcout(\Lab_UT.scdp.u0.byteToDecrypt_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22621),
            .ce(),
            .sr(N__18051));
    defparam \Lab_UT.scdp.u0.q_3_LC_5_14_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_3_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u0.q_3_LC_5_14_3 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \Lab_UT.scdp.u0.q_3_LC_5_14_3  (
            .in0(N__12952),
            .in1(N__11149),
            .in2(_gnd_net_),
            .in3(N__11161),
            .lcout(\Lab_UT.scdp.u0.byteToDecrypt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22621),
            .ce(),
            .sr(N__18051));
    defparam \Lab_UT.scdp.rxdataD.q_3_LC_5_14_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.rxdataD.q_3_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.rxdataD.q_3_LC_5_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.scdp.rxdataD.q_3_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11147),
            .lcout(\Lab_UT.scdp.binValD_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22621),
            .ce(),
            .sr(N__18051));
    defparam \Lab_UT.scdp.k1h.q_3_LC_5_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1h.q_3_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1h.q_3_LC_5_14_6 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.scdp.k1h.q_3_LC_5_14_6  (
            .in0(N__11121),
            .in1(N__15317),
            .in2(N__15249),
            .in3(N__13637),
            .lcout(\Lab_UT.scdp.key1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22621),
            .ce(),
            .sr(N__18051));
    defparam \Lab_UT.scdp.k1l.q_3_LC_5_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1l.q_3_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1l.q_3_LC_5_14_7 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \Lab_UT.scdp.k1l.q_3_LC_5_14_7  (
            .in0(N__15316),
            .in1(N__11106),
            .in2(N__15250),
            .in3(N__14200),
            .lcout(\Lab_UT.scdp.key1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22621),
            .ce(),
            .sr(N__18051));
    defparam \ufifo.txDataValidD_LC_5_15_0 .C_ON=1'b0;
    defparam \ufifo.txDataValidD_LC_5_15_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.txDataValidD_LC_5_15_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ufifo.txDataValidD_LC_5_15_0  (
            .in0(N__12661),
            .in1(N__12634),
            .in2(_gnd_net_),
            .in3(N__12655),
            .lcout(\ufifo.txDataValidDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22618),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIHLIO_3_LC_6_4_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIHLIO_3_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIHLIO_3_LC_6_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIHLIO_3_LC_6_4_1  (
            .in0(N__18309),
            .in1(N__20155),
            .in2(_gnd_net_),
            .in3(N__20095),
            .lcout(\Lab_UT.scctrl.g0_14_mb_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNI226B9_4_LC_6_5_0 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNI226B9_4_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNI226B9_4_LC_6_5_0 .LUT_INIT=16'b1110111011100000;
    LogicCell40 \ufifo.tx_fsm.cstate_RNI226B9_4_LC_6_5_0  (
            .in0(N__11225),
            .in1(N__11484),
            .in2(N__11523),
            .in3(N__21011),
            .lcout(),
            .ltout(\ufifo.N_57_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_1_LC_6_5_1 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_1_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \ufifo.emitcrlf_fsm.cstate_1_LC_6_5_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_1_LC_6_5_1  (
            .in0(N__11050),
            .in1(_gnd_net_),
            .in2(N__11044),
            .in3(N__11326),
            .lcout(\ufifo.emitcrlf_fsm.cstateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22661),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNI7ELR5_4_LC_6_5_2 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNI7ELR5_4_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNI7ELR5_4_LC_6_5_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ufifo.tx_fsm.cstate_RNI7ELR5_4_LC_6_5_2  (
            .in0(N__11513),
            .in1(N__11442),
            .in2(_gnd_net_),
            .in3(N__16184),
            .lcout(\ufifo.tx_fsm.N_59_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.shifter_ret_3_RNIP72B1_LC_6_5_3 .C_ON=1'b0;
    defparam \Lab_UT.dk.shifter_ret_3_RNIP72B1_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.shifter_ret_3_RNIP72B1_LC_6_5_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dk.shifter_ret_3_RNIP72B1_LC_6_5_3  (
            .in0(N__16297),
            .in1(N__16358),
            .in2(N__16171),
            .in3(N__16956),
            .lcout(\Lab_UT.m61_i_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.g0_LC_6_5_4 .C_ON=1'b0;
    defparam \Lab_UT.dk.g0_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.g0_LC_6_5_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dk.g0_LC_6_5_4  (
            .in0(N__11200),
            .in1(N__16162),
            .in2(_gnd_net_),
            .in3(N__20807),
            .lcout(\Lab_UT.de_bigE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_0_1_LC_6_5_5 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_0_1_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_0_1_LC_6_5_5 .LUT_INIT=16'b0101001100000000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNO_0_1_LC_6_5_5  (
            .in0(N__11443),
            .in1(N__12180),
            .in2(N__11385),
            .in3(N__20163),
            .lcout(\ufifo.emitcrlf_fsm.cstate_srsts_rn_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNO_0_0_LC_6_5_6 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNO_0_0_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNO_0_0_LC_6_5_6 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \ufifo.tx_fsm.cstate_RNO_0_0_LC_6_5_6  (
            .in0(N__11226),
            .in1(N__16185),
            .in2(_gnd_net_),
            .in3(N__21012),
            .lcout(),
            .ltout(\ufifo.tx_fsm.N_72_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_0_LC_6_5_7 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_0_LC_6_5_7 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_0_LC_6_5_7 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \ufifo.tx_fsm.cstate_0_LC_6_5_7  (
            .in0(N__11320),
            .in1(N__11302),
            .in2(N__11272),
            .in3(N__20164),
            .lcout(\ufifo.cstate_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22661),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNI6VBB5_LC_6_6_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNI6VBB5_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNI6VBB5_LC_6_6_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep2_RNI6VBB5_LC_6_6_0  (
            .in0(N__22305),
            .in1(N__20562),
            .in2(N__22093),
            .in3(N__17154),
            .lcout(\Lab_UT.scctrl.next_state_1_i_a5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.de_bigE_2_LC_6_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigE_2_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigE_2_LC_6_6_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dk.de_bigE_2_LC_6_6_1  (
            .in0(N__16510),
            .in1(N__16447),
            .in2(N__16971),
            .in3(N__17072),
            .lcout(\Lab_UT.dk.de_bigEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_6_6_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_6_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_6_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_18_LC_6_6_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_18_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_18_LC_6_6_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_18_LC_6_6_3  (
            .in0(N__14368),
            .in1(N__14433),
            .in2(_gnd_net_),
            .in3(N__20060),
            .lcout(\Lab_UT.scctrl.g0_i_a7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.state_ret_5_rep2_LC_6_6_6 .C_ON=1'b0;
    defparam \resetGen.state_ret_5_rep2_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \resetGen.state_ret_5_rep2_LC_6_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \resetGen.state_ret_5_rep2_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22762),
            .lcout(rst_i_3_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22654),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIMU571_2_LC_6_6_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIMU571_2_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIMU571_2_LC_6_6_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIMU571_2_LC_6_6_7  (
            .in0(N__20563),
            .in1(N__23001),
            .in2(N__19561),
            .in3(N__17502),
            .lcout(\Lab_UT.scctrl.un6_sccDecrypt ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_2_0_LC_6_7_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_2_0_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_2_0_LC_6_7_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_2_0_LC_6_7_0  (
            .in0(N__20786),
            .in1(N__11545),
            .in2(N__11641),
            .in3(N__13017),
            .lcout(\Lab_UT.scctrl.N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.de_cr_0_LC_6_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_cr_0_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_cr_0_LC_6_7_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dk.de_cr_0_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__16959),
            .in2(_gnd_net_),
            .in3(N__17066),
            .lcout(),
            .ltout(\Lab_UT.dk.escKey_4_reti_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.shifter_ret_3_LC_6_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dk.shifter_ret_3_LC_6_7_3 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dk.shifter_ret_3_LC_6_7_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \Lab_UT.dk.shifter_ret_3_LC_6_7_3  (
            .in0(N__13433),
            .in1(_gnd_net_),
            .in2(N__11539),
            .in3(N__15665),
            .lcout(\Lab_UT.de_cr_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22650),
            .ce(N__16757),
            .sr(N__18077));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_17_LC_6_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_17_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_17_LC_6_7_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_17_LC_6_7_4  (
            .in0(N__16353),
            .in1(N__16958),
            .in2(N__16292),
            .in3(N__16548),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_i_a3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_14_LC_6_7_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_14_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_14_LC_6_7_5 .LUT_INIT=16'b1100010001000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_14_LC_6_7_5  (
            .in0(N__22302),
            .in1(N__11536),
            .in2(N__11527),
            .in3(N__20785),
            .lcout(\Lab_UT.scctrl.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_a9_1_3_LC_6_7_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_a9_1_3_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_a9_1_3_LC_6_7_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_a9_1_3_LC_6_7_6  (
            .in0(N__16352),
            .in1(N__16155),
            .in2(N__16293),
            .in3(N__16957),
            .lcout(),
            .ltout(\Lab_UT.g0_i_a9_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_RNIQKK14_LC_6_7_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_RNIQKK14_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_11_RNIQKK14_LC_6_7_7 .LUT_INIT=16'b1100010001000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_RNIQKK14_LC_6_7_7  (
            .in0(N__22303),
            .in1(N__16060),
            .in2(N__11548),
            .in3(N__20784),
            .lcout(\Lab_UT.scctrl.N_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.shifter_ret_LC_6_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dk.shifter_ret_LC_6_8_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.dk.shifter_ret_LC_6_8_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \Lab_UT.dk.shifter_ret_LC_6_8_0  (
            .in0(N__13374),
            .in1(N__11897),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.de_cr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22644),
            .ce(N__16756),
            .sr(N__18073));
    defparam \buart.Z_rx.shifter_0_3_LC_6_8_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_3_LC_6_8_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_3_LC_6_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_3_LC_6_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13373),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22644),
            .ce(N__16756),
            .sr(N__18073));
    defparam \buart.Z_rx.shifter_0_fast_3_LC_6_8_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_3_LC_6_8_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_3_LC_6_8_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_fast_3_LC_6_8_2  (
            .in0(N__13375),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buart__rx_shifter_0_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22644),
            .ce(N__16756),
            .sr(N__18073));
    defparam \buart.Z_rx.shifter_0_0_LC_6_8_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_0_LC_6_8_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_0_LC_6_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_0_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15752),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22644),
            .ce(N__16756),
            .sr(N__18073));
    defparam \buart.Z_rx.shifter_0_1_LC_6_8_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_1_LC_6_8_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_1_LC_6_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_1_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15652),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22644),
            .ce(N__16756),
            .sr(N__18073));
    defparam \buart.Z_rx.shifter_0_0_rep1_LC_6_8_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_0_rep1_LC_6_8_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_0_rep1_LC_6_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_0_rep1_LC_6_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15753),
            .lcout(bu_rx_data_0_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22644),
            .ce(N__16756),
            .sr(N__18073));
    defparam \buart.Z_rx.shifter_ret_2_LC_6_8_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_2_LC_6_8_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_2_LC_6_8_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \buart.Z_rx.shifter_ret_2_LC_6_8_6  (
            .in0(_gnd_net_),
            .in1(N__16954),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22644),
            .ce(N__16756),
            .sr(N__18073));
    defparam \buart.Z_rx.shifter_0_2_LC_6_8_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_2_LC_6_8_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_2_LC_6_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_2_LC_6_8_7  (
            .in0(N__11898),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22644),
            .ce(N__16756),
            .sr(N__18073));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_2_LC_6_9_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_2_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_2_LC_6_9_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_2_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__12419),
            .in2(_gnd_net_),
            .in3(N__12372),
            .lcout(bu_rx_data_rdy),
            .ltout(bu_rx_data_rdy_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.r1.q_0_LC_6_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.r1.q_0_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.r1.q_0_LC_6_9_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \Lab_UT.scctrl.r1.q_0_LC_6_9_1  (
            .in0(N__17810),
            .in1(N__11569),
            .in2(N__11608),
            .in3(N__11563),
            .lcout(\Lab_UT.scctrl.delay1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22638),
            .ce(),
            .sr(N__18041));
    defparam \Lab_UT.scdp.pinst1.un1_pValid_LC_6_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.pinst1.un1_pValid_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.pinst1.un1_pValid_LC_6_9_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.scdp.pinst1.un1_pValid_LC_6_9_2  (
            .in0(N__13412),
            .in1(N__13305),
            .in2(_gnd_net_),
            .in3(N__16877),
            .lcout(\Lab_UT.un1_pValid ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.r2.q_0_LC_6_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.r2.q_0_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.r2.q_0_LC_6_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scctrl.r2.q_0_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11605),
            .lcout(\Lab_UT.scctrl.delay2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22638),
            .ce(),
            .sr(N__18041));
    defparam \Lab_UT.scctrl.r3.q_0_LC_6_9_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.r3.q_0_LC_6_9_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.r3.q_0_LC_6_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scctrl.r3.q_0_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11599),
            .lcout(\Lab_UT.scctrl.delay3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22638),
            .ce(),
            .sr(N__18041));
    defparam \Lab_UT.scdp.pinst1.un12_pValid_1_LC_6_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.pinst1.un12_pValid_1_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.pinst1.un12_pValid_1_LC_6_9_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scdp.pinst1.un12_pValid_1_LC_6_9_5  (
            .in0(N__13357),
            .in1(N__16354),
            .in2(_gnd_net_),
            .in3(N__13411),
            .lcout(),
            .ltout(\Lab_UT.scdp.pinst1.un12_pValidZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.pinst1.un7_pValid_LC_6_9_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.pinst1.un7_pValid_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.pinst1.un7_pValid_LC_6_9_6 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \Lab_UT.scdp.pinst1.un7_pValid_LC_6_9_6  (
            .in0(N__11586),
            .in1(N__16878),
            .in2(N__11572),
            .in3(N__17059),
            .lcout(\Lab_UT.un7_pValid ),
            .ltout(\Lab_UT.un7_pValid_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNIRB726_LC_6_9_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNIRB726_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNIRB726_LC_6_9_7 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNIRB726_LC_6_9_7  (
            .in0(N__17809),
            .in1(N__11562),
            .in2(N__11554),
            .in3(N__20753),
            .lcout(\Lab_UT.sccEldByte ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_6_RNIFERUH_LC_6_10_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_6_RNIFERUH_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_6_RNIFERUH_LC_6_10_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_6_RNIFERUH_LC_6_10_0  (
            .in0(N__21249),
            .in1(N__11713),
            .in2(N__21208),
            .in3(N__13583),
            .lcout(),
            .ltout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_6_RNIL97G01_LC_6_10_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_6_RNIL97G01_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_6_RNIL97G01_LC_6_10_1 .LUT_INIT=16'b0001001100010000;
    LogicCell40 \Lab_UT.scctrl.state_ret_6_RNIL97G01_LC_6_10_1  (
            .in0(N__13584),
            .in1(N__18939),
            .in2(N__11551),
            .in3(N__12786),
            .lcout(\Lab_UT.state_ret_6_RNIL97G01_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_0_sqmuxa_4_0_LC_6_10_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_0_sqmuxa_4_0_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_0_sqmuxa_4_0_LC_6_10_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.scctrl.next_state_0_sqmuxa_4_0_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21013),
            .in3(N__20209),
            .lcout(\Lab_UT.scctrl.next_state_0_sqmuxa_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.de_bigD_6_LC_6_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigD_6_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigD_6_LC_6_10_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dk.de_bigD_6_LC_6_10_3  (
            .in0(N__13252),
            .in1(N__11665),
            .in2(N__13473),
            .in3(N__13509),
            .lcout(Lab_UT_dk_de_bigD_6),
            .ltout(Lab_UT_dk_de_bigD_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.de_bigE_LC_6_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_bigE_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_bigE_LC_6_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dk.de_bigE_LC_6_10_4  (
            .in0(N__16136),
            .in1(N__11707),
            .in2(N__11701),
            .in3(N__20719),
            .lcout(\Lab_UT.de_bigE ),
            .ltout(\Lab_UT.de_bigE_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_6_RNIJMNGE_LC_6_10_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_6_RNIJMNGE_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_6_RNIJMNGE_LC_6_10_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Lab_UT.scctrl.state_ret_6_RNIJMNGE_LC_6_10_5  (
            .in0(N__13528),
            .in1(N__17135),
            .in2(N__11698),
            .in3(N__17198),
            .lcout(\Lab_UT.scctrl.next_state_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.val_i_0_LC_6_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_i_0_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_i_0_LC_6_11_0 .LUT_INIT=16'b0000101111110010;
    LogicCell40 \Lab_UT.scdp.a2b.val_i_0_LC_6_11_0  (
            .in0(N__14867),
            .in1(N__15680),
            .in2(N__11689),
            .in3(N__16146),
            .lcout(\Lab_UT.scdp.N_39 ),
            .ltout(\Lab_UT.scdp.N_39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.rxdataD.q_0_LC_6_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.rxdataD.q_0_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.rxdataD.q_0_LC_6_11_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \Lab_UT.scdp.rxdataD.q_0_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11695),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scdp.binValD_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22628),
            .ce(),
            .sr(N__18046));
    defparam \Lab_UT.scdp.a2b.val_0_o2_3_LC_6_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_0_o2_3_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_0_o2_3_LC_6_11_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \Lab_UT.scdp.a2b.val_0_o2_3_LC_6_11_2  (
            .in0(N__16879),
            .in1(N__13469),
            .in2(N__13324),
            .in3(N__11679),
            .lcout(\Lab_UT.scdp.a2b.N_50 ),
            .ltout(\Lab_UT.scdp.a2b.N_50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.val_i_o2_0_LC_6_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_i_o2_0_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_i_o2_0_LC_6_11_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.scdp.a2b.val_i_o2_0_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11692),
            .in3(N__11932),
            .lcout(\Lab_UT.scdp.a2b.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_8_0_LC_6_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_8_0_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_8_0_LC_6_11_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_8_0_LC_6_11_4  (
            .in0(N__14866),
            .in1(N__13468),
            .in2(N__11935),
            .in3(N__11678),
            .lcout(\Lab_UT.scctrl.m24_e_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.val_i_o2_1_LC_6_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_i_o2_1_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_i_o2_1_LC_6_11_5 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \Lab_UT.scdp.a2b.val_i_o2_1_LC_6_11_5  (
            .in0(N__11619),
            .in1(N__11933),
            .in2(_gnd_net_),
            .in3(N__16142),
            .lcout(\Lab_UT.scdp.a2b.N_53 ),
            .ltout(\Lab_UT.scdp.a2b.N_53_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.val_i_1_LC_6_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_i_1_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_i_1_LC_6_11_6 .LUT_INIT=16'b1010000010101100;
    LogicCell40 \Lab_UT.scdp.a2b.val_i_1_LC_6_11_6  (
            .in0(N__14868),
            .in1(N__15758),
            .in2(N__11872),
            .in3(N__15681),
            .lcout(\Lab_UT.scdp.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_0_LC_6_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_0_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u0.q_0_LC_6_11_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \Lab_UT.scdp.u0.q_0_LC_6_11_7  (
            .in0(N__11865),
            .in1(N__11838),
            .in2(_gnd_net_),
            .in3(N__12945),
            .lcout(\Lab_UT.scdp.byteToDecrypt_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22628),
            .ce(),
            .sr(N__18046));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_6_LC_6_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_6_LC_6_12_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_6_LC_6_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_6_LC_6_12_0  (
            .in0(N__11742),
            .in1(N__15529),
            .in2(_gnd_net_),
            .in3(N__12751),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22624),
            .ce(N__12467),
            .sr(N__18083));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNO_0_0_LC_6_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNO_0_0_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNO_0_0_LC_6_12_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNO_0_0_LC_6_12_1  (
            .in0(N__12500),
            .in1(N__11741),
            .in2(N__11823),
            .in3(N__11777),
            .lcout(),
            .ltout(\Lab_UT.scdp.lfsrInst.prng_lfsr_next_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_0_LC_6_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_0_LC_6_12_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_0_LC_6_12_2 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_0_LC_6_12_2  (
            .in0(N__13680),
            .in1(N__11796),
            .in2(N__11782),
            .in3(N__12748),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22624),
            .ce(N__12467),
            .sr(N__18083));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_2_LC_6_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_2_LC_6_12_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_2_LC_6_12_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_2_LC_6_12_3  (
            .in0(N__12747),
            .in1(N__13665),
            .in2(_gnd_net_),
            .in3(N__12522),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22624),
            .ce(N__12467),
            .sr(N__18083));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_5_LC_6_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_5_LC_6_12_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_5_LC_6_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_5_LC_6_12_4  (
            .in0(N__15838),
            .in1(N__11757),
            .in2(_gnd_net_),
            .in3(N__12750),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22624),
            .ce(N__12467),
            .sr(N__18083));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_12_LC_6_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_12_LC_6_12_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_12_LC_6_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_12_LC_6_12_5  (
            .in0(N__12745),
            .in1(N__13654),
            .in2(_gnd_net_),
            .in3(N__11725),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22624),
            .ce(N__12467),
            .sr(N__18083));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_1_LC_6_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_1_LC_6_12_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_1_LC_6_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_1_LC_6_12_6  (
            .in0(N__15343),
            .in1(N__12540),
            .in2(_gnd_net_),
            .in3(N__12749),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22624),
            .ce(N__12467),
            .sr(N__18083));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_13_LC_6_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_13_LC_6_12_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_13_LC_6_12_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_13_LC_6_12_7  (
            .in0(N__12746),
            .in1(_gnd_net_),
            .in2(N__12507),
            .in3(N__12613),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22624),
            .ce(N__12467),
            .sr(N__18083));
    defparam \Lab_UT.scdp.k3l.q_0_LC_6_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3l.q_0_LC_6_13_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3l.q_0_LC_6_13_0 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \Lab_UT.scdp.k3l.q_0_LC_6_13_0  (
            .in0(N__15497),
            .in1(N__12451),
            .in2(N__15272),
            .in3(N__13722),
            .lcout(\Lab_UT.scdp.key3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(),
            .sr(N__18052));
    defparam \Lab_UT.scdp.rddataDV.q_0_LC_6_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.rddataDV.q_0_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.rddataDV.q_0_LC_6_13_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.scdp.rddataDV.q_0_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(N__12439),
            .in2(_gnd_net_),
            .in3(N__12379),
            .lcout(\Lab_UT.scdp.binVal_ValidD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(),
            .sr(N__18052));
    defparam \Lab_UT.scdp.lsBitsi.q_0_LC_6_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_0_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_0_LC_6_13_2 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_0_LC_6_13_2  (
            .in0(N__13181),
            .in1(N__12361),
            .in2(N__12333),
            .in3(N__12313),
            .lcout(\Lab_UT.scdp.lsBitsD_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(),
            .sr(N__18052));
    defparam \Lab_UT.scdp.lsBitsi.q_4_LC_6_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_4_LC_6_13_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_4_LC_6_13_3 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_4_LC_6_13_3  (
            .in0(N__12285),
            .in1(N__12312),
            .in2(_gnd_net_),
            .in3(N__13183),
            .lcout(\Lab_UT.scdp.lsBitsD_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(),
            .sr(N__18052));
    defparam \Lab_UT.scdp.msBitsi.q_3_LC_6_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_3_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_3_LC_6_13_4 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_3_LC_6_13_4  (
            .in0(N__13182),
            .in1(N__12268),
            .in2(N__12207),
            .in3(N__12229),
            .lcout(\Lab_UT.scdp.msBitsD_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(),
            .sr(N__18052));
    defparam \buart.Z_tx.bitcount_0_LC_6_13_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_6_13_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_6_13_5 .LUT_INIT=16'b0110101000000000;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_6_13_5  (
            .in0(N__11960),
            .in1(N__12184),
            .in2(N__12115),
            .in3(N__12052),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(),
            .sr(N__18052));
    defparam \Lab_UT.scctrl.state_ret_13_RNIQ72741_LC_6_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNIQ72741_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNIQ72741_LC_6_13_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNIQ72741_LC_6_13_6  (
            .in0(N__13638),
            .in1(N__15034),
            .in2(_gnd_net_),
            .in3(N__14983),
            .lcout(\Lab_UT.state_ret_13_RNIQ72741_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.r4.q_0_LC_6_13_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.r4.q_0_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.r4.q_0_LC_6_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scctrl.r4.q_0_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12654),
            .lcout(\Lab_UT.scctrl.r4.delay4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(),
            .sr(N__18052));
    defparam \Lab_UT.scdp.u1.q_esr_2_LC_6_14_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_esr_2_LC_6_14_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u1.q_esr_2_LC_6_14_0 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \Lab_UT.scdp.u1.q_esr_2_LC_6_14_0  (
            .in0(N__15682),
            .in1(N__15776),
            .in2(_gnd_net_),
            .in3(N__15809),
            .lcout(\Lab_UT.scdp.u1.byteToDecrypt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22617),
            .ce(N__14047),
            .sr(N__18054));
    defparam \Lab_UT.scctrl.state_2_RNI44QH41_2_LC_6_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNI44QH41_2_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNI44QH41_2_LC_6_14_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scctrl.state_2_RNI44QH41_2_LC_6_14_5  (
            .in0(N__13771),
            .in1(N__18199),
            .in2(_gnd_net_),
            .in3(N__14984),
            .lcout(\Lab_UT.state_2_RNI44QH41_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNI416G41_LC_6_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNI416G41_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNI416G41_LC_6_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNI416G41_LC_6_14_6  (
            .in0(N__14986),
            .in1(N__14676),
            .in2(_gnd_net_),
            .in3(N__13837),
            .lcout(\Lab_UT.state_ret_14_RNI416G41_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIF0RJ41_2_LC_6_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIF0RJ41_2_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIF0RJ41_2_LC_6_14_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIF0RJ41_2_LC_6_14_7  (
            .in0(N__13726),
            .in1(N__18220),
            .in2(_gnd_net_),
            .in3(N__14985),
            .lcout(\Lab_UT.state_2_RNIF0RJ41_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.k1h.q_1_LC_6_15_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1h.q_1_LC_6_15_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1h.q_1_LC_6_15_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.scdp.k1h.q_1_LC_6_15_0  (
            .in0(N__12612),
            .in1(N__15384),
            .in2(N__15274),
            .in3(N__13639),
            .lcout(\Lab_UT.scdp.key1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22615),
            .ce(),
            .sr(N__18055));
    defparam \Lab_UT.scdp.k1l.q_1_LC_6_15_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1l.q_1_LC_6_15_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1l.q_1_LC_6_15_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.scdp.k1l.q_1_LC_6_15_1  (
            .in0(N__15383),
            .in1(N__15231),
            .in2(N__12597),
            .in3(N__14199),
            .lcout(\Lab_UT.scdp.key1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22615),
            .ce(),
            .sr(N__18055));
    defparam \Lab_UT.scdp.k2h.q_1_LC_6_15_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2h.q_1_LC_6_15_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2h.q_1_LC_6_15_2 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.scdp.k2h.q_1_LC_6_15_2  (
            .in0(N__12573),
            .in1(N__15385),
            .in2(N__15275),
            .in3(N__13768),
            .lcout(\Lab_UT.scdp.key2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22615),
            .ce(),
            .sr(N__18055));
    defparam \Lab_UT.scdp.k3h.q_1_LC_6_15_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3h.q_1_LC_6_15_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3h.q_1_LC_6_15_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \Lab_UT.scdp.k3h.q_1_LC_6_15_3  (
            .in0(N__13835),
            .in1(N__15233),
            .in2(N__15391),
            .in3(N__12558),
            .lcout(\Lab_UT.scdp.key3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22615),
            .ce(),
            .sr(N__18055));
    defparam \Lab_UT.scdp.k3l.q_1_LC_6_15_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3l.q_1_LC_6_15_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3l.q_1_LC_6_15_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k3l.q_1_LC_6_15_4  (
            .in0(N__15229),
            .in1(N__15386),
            .in2(N__12906),
            .in3(N__13723),
            .lcout(\Lab_UT.scdp.key3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22615),
            .ce(),
            .sr(N__18055));
    defparam \Lab_UT.scdp.k1l.q_0_LC_6_15_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1l.q_0_LC_6_15_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1l.q_0_LC_6_15_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.scdp.k1l.q_0_LC_6_15_5  (
            .in0(N__15498),
            .in1(N__15230),
            .in2(N__12885),
            .in3(N__14198),
            .lcout(\Lab_UT.scdp.key1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22615),
            .ce(),
            .sr(N__18055));
    defparam \Lab_UT.scdp.k2h.q_0_LC_6_15_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2h.q_0_LC_6_15_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2h.q_0_LC_6_15_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k2h.q_0_LC_6_15_6  (
            .in0(N__15228),
            .in1(N__15499),
            .in2(N__12865),
            .in3(N__13767),
            .lcout(\Lab_UT.scdp.key2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22615),
            .ce(),
            .sr(N__18055));
    defparam \Lab_UT.scdp.k3h.q_0_LC_6_15_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3h.q_0_LC_6_15_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3h.q_0_LC_6_15_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \Lab_UT.scdp.k3h.q_0_LC_6_15_7  (
            .in0(N__13834),
            .in1(N__15232),
            .in2(N__15509),
            .in3(N__12837),
            .lcout(\Lab_UT.scdp.key3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22615),
            .ce(),
            .sr(N__18055));
    defparam \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_LC_6_16_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_LC_6_16_0 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_LC_6_16_0  (
            .in0(N__12819),
            .in1(N__14117),
            .in2(N__14155),
            .in3(N__12744),
            .lcout(\Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNIMEE3_LC_6_16_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNIMEE3_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNIMEE3_LC_6_16_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNIMEE3_LC_6_16_2  (
            .in0(N__22268),
            .in1(N__19698),
            .in2(_gnd_net_),
            .in3(N__21955),
            .lcout(),
            .ltout(\Lab_UT.scctrl.un1_state_inv_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_12_RNIUQFK_LC_6_16_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_12_RNIUQFK_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_12_RNIUQFK_LC_6_16_3 .LUT_INIT=16'b0111111101110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_12_RNIUQFK_LC_6_16_3  (
            .in0(N__20256),
            .in1(N__20577),
            .in2(N__12670),
            .in3(N__18955),
            .lcout(),
            .ltout(\Lab_UT.scctrl.state_ret_12_RNIUQFKZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_12_RNIMJCP8_LC_6_16_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_12_RNIMJCP8_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_12_RNIMJCP8_LC_6_16_4 .LUT_INIT=16'b0000110000001110;
    LogicCell40 \Lab_UT.scctrl.state_ret_12_RNIMJCP8_LC_6_16_4  (
            .in0(N__13048),
            .in1(N__14118),
            .in2(N__12667),
            .in3(N__19150),
            .lcout(\Lab_UT.state_ret_12_RNIMJCP8_0 ),
            .ltout(\Lab_UT.state_ret_12_RNIMJCP8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.r5.q_0_LC_6_16_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.r5.q_0_LC_6_16_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.r5.q_0_LC_6_16_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \Lab_UT.scctrl.r5.q_0_LC_6_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12664),
            .in3(N__14153),
            .lcout(\Lab_UT.scctrl.delayload ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22614),
            .ce(),
            .sr(N__18058));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_5_LC_6_16_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_5_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_5_LC_6_16_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_5_LC_6_16_7  (
            .in0(N__19699),
            .in1(N__20576),
            .in2(_gnd_net_),
            .in3(N__22269),
            .lcout(\Lab_UT.scctrl.g0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNIM6P13_LC_7_3_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNIM6P13_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNIM6P13_LC_7_3_1 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNIM6P13_LC_7_3_1  (
            .in0(N__21127),
            .in1(N__17623),
            .in2(_gnd_net_),
            .in3(N__21014),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNISBDB3_2_LC_7_3_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNISBDB3_2_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNISBDB3_2_LC_7_3_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.scctrl.next_state_RNISBDB3_2_LC_7_3_2  (
            .in0(N__20084),
            .in1(_gnd_net_),
            .in2(N__12922),
            .in3(N__20308),
            .lcout(\Lab_UT.scctrl.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNINMBN3_LC_7_3_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNINMBN3_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNINMBN3_LC_7_3_4 .LUT_INIT=16'b1000000010001000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNINMBN3_LC_7_3_4  (
            .in0(N__20083),
            .in1(N__19695),
            .in2(N__13495),
            .in3(N__20803),
            .lcout(\Lab_UT.scctrl.g0_i_a9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNI07T4_LC_7_3_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNI07T4_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNI07T4_LC_7_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNI07T4_LC_7_3_5  (
            .in0(N__19696),
            .in1(N__20082),
            .in2(N__22339),
            .in3(N__20462),
            .lcout(\Lab_UT.scctrl.G_23_0_a9_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNI4DGV4_LC_7_3_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNI4DGV4_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNI4DGV4_LC_7_3_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNI4DGV4_LC_7_3_6  (
            .in0(N__14206),
            .in1(N__13552),
            .in2(N__16408),
            .in3(N__20804),
            .lcout(\Lab_UT.scctrl.g0_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.state_ret_5_rep1_LC_7_4_2 .C_ON=1'b0;
    defparam \resetGen.state_ret_5_rep1_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.state_ret_5_rep1_LC_7_4_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \resetGen.state_ret_5_rep1_LC_7_4_2  (
            .in0(N__22768),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rst_i_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22679),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIO386G1_2_LC_7_4_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIO386G1_2_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIO386G1_2_LC_7_4_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIO386G1_2_LC_7_4_3  (
            .in0(N__14473),
            .in1(N__14346),
            .in2(_gnd_net_),
            .in3(N__14331),
            .lcout(),
            .ltout(\Lab_UT.scctrl.un1_state_3_1_reti_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_10_LC_7_4_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_10_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_10_LC_7_4_4 .LUT_INIT=16'b0111010101010101;
    LogicCell40 \Lab_UT.scctrl.state_ret_10_LC_7_4_4  (
            .in0(N__22767),
            .in1(N__14212),
            .in2(N__12919),
            .in3(N__14290),
            .lcout(\Lab_UT.scctrl.state_retZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22679),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNI0D9CA_LC_7_4_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNI0D9CA_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNI0D9CA_LC_7_4_5 .LUT_INIT=16'b0100000001000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNI0D9CA_LC_7_4_5  (
            .in0(N__18947),
            .in1(N__20076),
            .in2(N__12916),
            .in3(N__13021),
            .lcout(\Lab_UT.scctrl.g0_16_mb_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.state_ret_5_LC_7_5_0 .C_ON=1'b0;
    defparam \resetGen.state_ret_5_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.state_ret_5_LC_7_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \resetGen.state_ret_5_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22780),
            .lcout(rst_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22674),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_11_LC_7_5_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_11_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_11_LC_7_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_11_LC_7_5_1  (
            .in0(N__21424),
            .in1(N__20075),
            .in2(N__21782),
            .in3(N__22090),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_4_LC_7_5_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_4_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_4_LC_7_5_2 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_4_LC_7_5_2  (
            .in0(N__12994),
            .in1(N__19425),
            .in2(N__12985),
            .in3(N__21006),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_1_LC_7_5_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_1_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_1_LC_7_5_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_1_LC_7_5_3  (
            .in0(N__12961),
            .in1(N__12976),
            .in2(N__12982),
            .in3(N__18967),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_0_LC_7_5_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_0_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_0_LC_7_5_4 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_0_LC_7_5_4  (
            .in0(N__12970),
            .in1(N__14289),
            .in2(N__12979),
            .in3(N__14521),
            .lcout(\Lab_UT.scctrl.N_1_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_6_LC_7_5_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_6_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_6_LC_7_5_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_6_LC_7_5_5  (
            .in0(N__20077),
            .in1(N__23021),
            .in2(N__21439),
            .in3(N__19166),
            .lcout(\Lab_UT.scctrl.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_2_LC_7_5_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_2_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_2_LC_7_5_6 .LUT_INIT=16'b0000001111110011;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_2_LC_7_5_6  (
            .in0(_gnd_net_),
            .in1(N__20331),
            .in2(N__20097),
            .in3(N__17888),
            .lcout(\Lab_UT.scctrl.g2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_7_LC_7_5_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_7_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_7_LC_7_5_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_7_LC_7_5_7  (
            .in0(N__21007),
            .in1(_gnd_net_),
            .in2(N__21173),
            .in3(N__20071),
            .lcout(\Lab_UT.scctrl.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_10_RNIPCFBB_LC_7_6_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_10_RNIPCFBB_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_10_RNIPCFBB_LC_7_6_0 .LUT_INIT=16'b0010001100000001;
    LogicCell40 \Lab_UT.scctrl.state_ret_10_RNIPCFBB_LC_7_6_0  (
            .in0(N__13110),
            .in1(N__14146),
            .in2(N__13096),
            .in3(N__13059),
            .lcout(\Lab_UT.sccDnibble1En ),
            .ltout(\Lab_UT.sccDnibble1En_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_esr_RNO_2_LC_7_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_esr_RNO_2_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_esr_RNO_2_LC_7_6_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.scdp.u0.q_esr_RNO_2_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13129),
            .in3(N__14087),
            .lcout(\Lab_UT.scdp.u0.sccDnibble1En_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_RNI658G_LC_7_6_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNI658G_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNI658G_LC_7_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNI658G_LC_7_6_2  (
            .in0(N__21742),
            .in1(N__17554),
            .in2(N__21440),
            .in3(N__21927),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_1_sqmuxa_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_RNI4CFD9_LC_7_6_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNI4CFD9_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNI4CFD9_LC_7_6_3 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNI4CFD9_LC_7_6_3  (
            .in0(N__18612),
            .in1(_gnd_net_),
            .in2(N__13114),
            .in3(N__18771),
            .lcout(\Lab_UT.scctrl.next_state_1_sqmuxa_3 ),
            .ltout(\Lab_UT.scctrl.next_state_1_sqmuxa_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_LC_7_6_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_LC_7_6_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.nibbleIn1_LC_7_6_4 .LUT_INIT=16'b0111111100001000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_LC_7_6_4  (
            .in0(N__13111),
            .in1(N__22781),
            .in2(N__13099),
            .in3(N__13095),
            .lcout(\Lab_UT.scctrl.nibbleInZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22666),
            .ce(N__13081),
            .sr(N__13066));
    defparam \Lab_UT.scctrl.state_ret_8_RNIQ79K1_LC_7_6_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNIQ79K1_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNIQ79K1_LC_7_6_5 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNIQ79K1_LC_7_6_5  (
            .in0(N__13044),
            .in1(N__21950),
            .in2(N__21791),
            .in3(N__21428),
            .lcout(\Lab_UT.sccDecrypt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_11_LC_7_6_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_11_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_11_LC_7_6_6 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_11_LC_7_6_6  (
            .in0(N__21743),
            .in1(N__18611),
            .in2(N__14278),
            .in3(N__18763),
            .lcout(\Lab_UT.scctrl.N_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_RNIJLL09_LC_7_6_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNIJLL09_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNIJLL09_LC_7_6_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNIJLL09_LC_7_6_7  (
            .in0(N__18764),
            .in1(N__15985),
            .in2(N__18627),
            .in3(N__21949),
            .lcout(\Lab_UT.scctrl.N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIHB2UD_LC_7_7_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIHB2UD_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIHB2UD_LC_7_7_0 .LUT_INIT=16'b0010101000111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNIHB2UD_LC_7_7_0  (
            .in0(N__13030),
            .in1(N__20928),
            .in2(N__14269),
            .in3(N__13016),
            .lcout(\Lab_UT.next_state_rst_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNIK9603_LC_7_7_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNIK9603_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNIK9603_LC_7_7_2 .LUT_INIT=16'b0101010100010000;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNIK9603_LC_7_7_2  (
            .in0(N__18913),
            .in1(N__20927),
            .in2(N__17840),
            .in3(N__13000),
            .lcout(\Lab_UT.scctrl.EmsLoaded ),
            .ltout(\Lab_UT.scctrl.EmsLoaded_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNIEOE1_LC_7_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNIEOE1_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNIEOE1_LC_7_7_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNIEOE1_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13210),
            .in3(N__17829),
            .lcout(\Lab_UT.sccElsBitsLd ),
            .ltout(\Lab_UT.sccElsBitsLd_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_ctle_6_LC_7_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_ctle_6_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_ctle_6_LC_7_7_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_ctle_6_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13207),
            .in3(N__14094),
            .lcout(\Lab_UT.scdp.sccElsBitsLd_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNO_6_LC_7_7_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_6_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_6_LC_7_7_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNO_6_LC_7_7_6  (
            .in0(N__18914),
            .in1(N__20184),
            .in2(_gnd_net_),
            .in3(N__20078),
            .lcout(\Lab_UT.scctrl.G_24_i_a4_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lsBitsi.q_5_LC_7_7_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_5_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_5_LC_7_7_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_5_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(N__13146),
            .in2(_gnd_net_),
            .in3(N__13170),
            .lcout(\Lab_UT.scdp.lsBitsi.lsBitsD_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22659),
            .ce(),
            .sr(N__18044));
    defparam \Lab_UT.dk.shifter_ret_3_RNIA82U_LC_7_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dk.shifter_ret_3_RNIA82U_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.shifter_ret_3_RNIA82U_LC_7_8_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dk.shifter_ret_3_RNIA82U_LC_7_8_0  (
            .in0(N__16270),
            .in1(N__16341),
            .in2(_gnd_net_),
            .in3(N__16944),
            .lcout(Lab_UT_dk_de_cr_12_1),
            .ltout(Lab_UT_dk_de_cr_12_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.shifter_ret_3_RNIJC3U2_LC_7_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dk.shifter_ret_3_RNIJC3U2_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.shifter_ret_3_RNIJC3U2_LC_7_8_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \Lab_UT.dk.shifter_ret_3_RNIJC3U2_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__16546),
            .in2(N__13135),
            .in3(N__20718),
            .lcout(L4_PrintBuf),
            .ltout(L4_PrintBuf_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIHA8U3_LC_7_8_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIHA8U3_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIHA8U3_LC_7_8_2 .LUT_INIT=16'b0101010111110101;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep1_RNIHA8U3_LC_7_8_2  (
            .in0(N__17576),
            .in1(_gnd_net_),
            .in2(N__13132),
            .in3(N__14701),
            .lcout(\Lab_UT.state_ret_8_rep1_RNIHA8U3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI5GLD_0_3_LC_7_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI5GLD_0_3_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI5GLD_0_3_LC_7_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI5GLD_0_3_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__20521),
            .in2(_gnd_net_),
            .in3(N__17499),
            .lcout(\Lab_UT.scctrl.g0_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.g1_i_a7_2_3_LC_7_8_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.g1_i_a7_2_3_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.g1_i_a7_2_3_LC_7_8_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.scctrl.g1_i_a7_2_3_LC_7_8_4  (
            .in0(N__16547),
            .in1(N__16342),
            .in2(N__16291),
            .in3(N__16945),
            .lcout(\Lab_UT.scctrl.g1_i_a7_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_8_LC_7_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_8_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_8_LC_7_8_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_8_LC_7_8_5  (
            .in0(N__20911),
            .in1(N__20018),
            .in2(N__21200),
            .in3(N__13264),
            .lcout(\Lab_UT.scctrl.g0_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI6J7KA_3_LC_7_8_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI6J7KA_3_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI6J7KA_3_LC_7_8_6 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI6J7KA_3_LC_7_8_6  (
            .in0(N__17500),
            .in1(N__19069),
            .in2(N__23073),
            .in3(N__20910),
            .lcout(\Lab_UT.N_190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g1_1_o2_0_0_LC_7_8_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g1_1_o2_0_0_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g1_1_o2_0_0_LC_7_8_7 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \Lab_UT.scdp.a2b.g1_1_o2_0_0_LC_7_8_7  (
            .in0(N__20912),
            .in1(N__14404),
            .in2(N__19118),
            .in3(N__13519),
            .lcout(\Lab_UT.scdp.a2b.g1_1_o2_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_fast_0_LC_7_9_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_0_LC_7_9_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_0_LC_7_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_fast_0_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15754),
            .lcout(bu_rx_data_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22647),
            .ce(N__16755),
            .sr(N__18079));
    defparam \Lab_UT.dk.un7_de_hex_x0_LC_7_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dk.un7_de_hex_x0_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.un7_de_hex_x0_LC_7_9_1 .LUT_INIT=16'b0000101000010011;
    LogicCell40 \Lab_UT.dk.un7_de_hex_x0_LC_7_9_1  (
            .in0(N__16500),
            .in1(N__13216),
            .in2(N__13510),
            .in3(N__13258),
            .lcout(),
            .ltout(\Lab_UT.dk.un7_de_hex_xZ0Z0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.un7_de_hex_ns_LC_7_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dk.un7_de_hex_ns_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.un7_de_hex_ns_LC_7_9_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.dk.un7_de_hex_ns_LC_7_9_2  (
            .in0(N__13251),
            .in1(_gnd_net_),
            .in2(N__13231),
            .in3(N__13964),
            .lcout(\Lab_UT.dk.un7_de_hex_0 ),
            .ltout(\Lab_UT.dk.un7_de_hex_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.de_hex_LC_7_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dk.de_hex_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.de_hex_LC_7_9_3 .LUT_INIT=16'b0111001101110111;
    LogicCell40 \Lab_UT.dk.de_hex_LC_7_9_3  (
            .in0(N__13278),
            .in1(N__20713),
            .in2(N__13228),
            .in3(N__13483),
            .lcout(\Lab_UT.de_hex_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.un4_de_hex_LC_7_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dk.un4_de_hex_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.un4_de_hex_LC_7_9_4 .LUT_INIT=16'b0010000000100000;
    LogicCell40 \Lab_UT.dk.un4_de_hex_LC_7_9_4  (
            .in0(N__13482),
            .in1(N__13225),
            .in2(N__20757),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.un4_de_hex ),
            .ltout(\Lab_UT.un4_de_hex_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNI68R1A_2_LC_7_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNI68R1A_2_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNI68R1A_2_LC_7_9_5 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNI68R1A_2_LC_7_9_5  (
            .in0(N__20752),
            .in1(N__14359),
            .in2(N__13219),
            .in3(N__13279),
            .lcout(\Lab_UT.N_191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_fast_1_LC_7_9_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_1_LC_7_9_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_1_LC_7_9_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_fast_1_LC_7_9_6  (
            .in0(N__15651),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buart__rx_shifter_0_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22647),
            .ce(N__16755),
            .sr(N__18079));
    defparam \buart.Z_rx.shifter_ret_1_fast_LC_7_9_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_1_fast_LC_7_9_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_1_fast_LC_7_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_1_fast_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15650),
            .lcout(buart__rx_shifter_ret_1_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22647),
            .ce(N__16755),
            .sr(N__18079));
    defparam \Lab_UT.scctrl.g0_i_o9_0_2_LC_7_10_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.g0_i_o9_0_2_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.g0_i_o9_0_2_LC_7_10_0 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \Lab_UT.scctrl.g0_i_o9_0_2_LC_7_10_0  (
            .in0(N__13408),
            .in1(N__13350),
            .in2(N__13323),
            .in3(N__16890),
            .lcout(\Lab_UT.scctrl.g0_i_o9_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_4_LC_7_10_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_4_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_4_LC_7_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_4_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13410),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22641),
            .ce(N__16758),
            .sr(N__18081));
    defparam \buart.Z_rx.shifter_0_5_LC_7_10_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_5_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_5_LC_7_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_5_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17049),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22641),
            .ce(N__16758),
            .sr(N__18081));
    defparam \Lab_UT.dk.un4_de_hex_1_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dk.un4_de_hex_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.un4_de_hex_1_LC_7_10_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dk.un4_de_hex_1_LC_7_10_3  (
            .in0(N__17048),
            .in1(N__13406),
            .in2(N__16940),
            .in3(N__13464),
            .lcout(\Lab_UT.dk.un4_de_hexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_ret_LC_7_10_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_LC_7_10_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_LC_7_10_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_LC_7_10_4  (
            .in0(N__13409),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22641),
            .ce(N__16758),
            .sr(N__18081));
    defparam \Lab_UT.dk.un1_de_hex_2_LC_7_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dk.un1_de_hex_2_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.un1_de_hex_2_LC_7_10_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dk.un1_de_hex_2_LC_7_10_6  (
            .in0(N__13407),
            .in1(N__13349),
            .in2(N__13322),
            .in3(N__16886),
            .lcout(\Lab_UT.un1_de_hex_2 ),
            .ltout(\Lab_UT.un1_de_hex_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.un1_de_hex_LC_7_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dk.un1_de_hex_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dk.un1_de_hex_LC_7_10_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.dk.un1_de_hex_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13267),
            .in3(N__20717),
            .lcout(\Lab_UT.un1_de_hex ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI55RL_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI55RL_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI55RL_LC_7_11_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_fast_RNI55RL_LC_7_11_0  (
            .in0(N__16941),
            .in1(N__19915),
            .in2(N__14443),
            .in3(N__19211),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_i_a9_3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI86TJ1_LC_7_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI86TJ1_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI86TJ1_LC_7_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_fast_RNI86TJ1_LC_7_11_1  (
            .in0(N__16164),
            .in1(N__16305),
            .in2(N__13555),
            .in3(N__16367),
            .lcout(\Lab_UT.scctrl.g0_i_a9_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNO_9_LC_7_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_9_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_9_LC_7_11_2 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNO_9_LC_7_11_2  (
            .in0(N__16942),
            .in1(N__16165),
            .in2(N__16372),
            .in3(N__16306),
            .lcout(\Lab_UT.scctrl.m26_i_o4_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI7JDJ_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI7JDJ_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI7JDJ_LC_7_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_fast_RNI7JDJ_LC_7_11_3  (
            .in0(N__19212),
            .in1(N__14442),
            .in2(_gnd_net_),
            .in3(N__21673),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_1_0_a5_2_out_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI21I2A_LC_7_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI21I2A_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_fast_RNI21I2A_LC_7_11_4 .LUT_INIT=16'b0000010100010101;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_fast_RNI21I2A_LC_7_11_4  (
            .in0(N__13915),
            .in1(N__18591),
            .in2(N__13537),
            .in3(N__18730),
            .lcout(\Lab_UT.next_state_1_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_0_1_LC_7_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_0_1_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_0_1_LC_7_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.scctrl.state_0_1_LC_7_11_5  (
            .in0(N__19916),
            .in1(N__17686),
            .in2(_gnd_net_),
            .in3(N__14622),
            .lcout(\Lab_UT.state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22635),
            .ce(),
            .sr(N__18048));
    defparam \Lab_UT.scctrl.state_ret_LC_7_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_LC_7_11_6 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_LC_7_11_6  (
            .in0(N__14623),
            .in1(N__17687),
            .in2(N__14482),
            .in3(N__19917),
            .lcout(\Lab_UT.scctrl.N_222_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22635),
            .ce(),
            .sr(N__18048));
    defparam \Lab_UT.scctrl.state_ret_RNILUJH_LC_7_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_RNILUJH_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_RNILUJH_LC_7_11_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_RNILUJH_LC_7_11_7  (
            .in0(N__19662),
            .in1(N__21941),
            .in2(_gnd_net_),
            .in3(N__13534),
            .lcout(\Lab_UT.scctrl.next_state76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_6_RNICI45_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_6_RNICI45_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_6_RNICI45_LC_7_12_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_6_RNICI45_LC_7_12_1  (
            .in0(N__21426),
            .in1(N__21248),
            .in2(_gnd_net_),
            .in3(N__17343),
            .lcout(\Lab_UT.scctrl.next_state_3_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g1_1_a3_0_0_LC_7_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g1_1_a3_0_0_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g1_1_a3_0_0_LC_7_12_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.scdp.a2b.g1_1_a3_0_0_LC_7_12_3  (
            .in0(N__21427),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23088),
            .lcout(\Lab_UT.scdp.a2b.g1_1_a3_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.k0l.q_0_LC_7_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0l.q_0_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0l.q_0_LC_7_12_4 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \Lab_UT.scdp.k0l.q_0_LC_7_12_4  (
            .in0(N__15489),
            .in1(N__13681),
            .in2(N__15276),
            .in3(N__15075),
            .lcout(\Lab_UT.scdp.key0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22630),
            .ce(),
            .sr(N__18053));
    defparam \Lab_UT.scdp.k0l.q_2_LC_7_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0l.q_2_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0l.q_2_LC_7_12_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.scdp.k0l.q_2_LC_7_12_5  (
            .in0(N__15076),
            .in1(N__15240),
            .in2(N__13669),
            .in3(N__15567),
            .lcout(\Lab_UT.scdp.key0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22630),
            .ce(),
            .sr(N__18053));
    defparam \Lab_UT.scdp.k1h.q_0_LC_7_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1h.q_0_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1h.q_0_LC_7_12_6 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \Lab_UT.scdp.k1h.q_0_LC_7_12_6  (
            .in0(N__15490),
            .in1(N__13653),
            .in2(N__15277),
            .in3(N__13636),
            .lcout(\Lab_UT.scdp.key1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22630),
            .ce(),
            .sr(N__18053));
    defparam \Lab_UT.scdp.k1h.q_2_LC_7_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1h.q_2_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1h.q_2_LC_7_12_7 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Lab_UT.scdp.k1h.q_2_LC_7_12_7  (
            .in0(N__13635),
            .in1(N__13602),
            .in2(N__15286),
            .in3(N__15568),
            .lcout(\Lab_UT.scdp.key1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22630),
            .ce(),
            .sr(N__18053));
    defparam \Lab_UT.scctrl.state_0_RNIBE791_1_LC_7_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_0_RNIBE791_1_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_0_RNIBE791_1_LC_7_13_0 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \Lab_UT.scctrl.state_0_RNIBE791_1_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__21698),
            .in2(N__23094),
            .in3(N__13911),
            .lcout(\Lab_UT.scctrl.next_state77 ),
            .ltout(\Lab_UT.scctrl.next_state77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_3_RNIHF1E3_LC_7_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_3_RNIHF1E3_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_3_RNIHF1E3_LC_7_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.scctrl.state_ret_3_RNIHF1E3_LC_7_13_1  (
            .in0(N__13884),
            .in1(N__14727),
            .in2(N__13588),
            .in3(N__14995),
            .lcout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNIG62DM_LC_7_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNIG62DM_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNIG62DM_LC_7_13_2 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNIG62DM_LC_7_13_2  (
            .in0(N__15030),
            .in1(N__19108),
            .in2(N__20222),
            .in3(N__13585),
            .lcout(),
            .ltout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNI91DN31_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNI91DN31_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNI91DN31_LC_7_13_3 .LUT_INIT=16'b0000111101001111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNI91DN31_LC_7_13_3  (
            .in0(N__19109),
            .in1(N__20188),
            .in2(N__13567),
            .in3(N__13894),
            .lcout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i ),
            .ltout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_0_RNIKFK051_1_LC_7_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_0_RNIKFK051_1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_0_RNIKFK051_1_LC_7_13_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \Lab_UT.scctrl.state_0_RNIKFK051_1_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__13564),
            .in2(N__13558),
            .in3(N__15081),
            .lcout(\Lab_UT.state_0_RNIKFK051_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep1_RNIT6TH_LC_7_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep1_RNIT6TH_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep1_RNIT6TH_LC_7_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep1_RNIT6TH_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__19210),
            .in2(_gnd_net_),
            .in3(N__17440),
            .lcout(\Lab_UT.scctrl.next_state77_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIDHLT5_2_LC_7_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIDHLT5_2_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIDHLT5_2_LC_7_13_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIDHLT5_2_LC_7_13_6  (
            .in0(N__18198),
            .in1(N__18216),
            .in2(N__14677),
            .in3(N__13900),
            .lcout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_RNIUV0941_LC_7_13_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_RNIUV0941_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_RNIUV0941_LC_7_13_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_RNIUV0941_LC_7_13_7  (
            .in0(N__15433),
            .in1(_gnd_net_),
            .in2(N__13888),
            .in3(N__14982),
            .lcout(\Lab_UT.state_ret_RNIUV0941_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.k2l.q_3_LC_7_14_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2l.q_3_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2l.q_3_LC_7_14_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.scdp.k2l.q_3_LC_7_14_0  (
            .in0(N__13869),
            .in1(N__15322),
            .in2(N__15251),
            .in3(N__14911),
            .lcout(\Lab_UT.scdp.key2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22622),
            .ce(),
            .sr(N__18056));
    defparam \Lab_UT.scdp.k2h.q_2_LC_7_14_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2h.q_2_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2h.q_2_LC_7_14_1 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.scdp.k2h.q_2_LC_7_14_1  (
            .in0(N__13851),
            .in1(N__15558),
            .in2(N__15247),
            .in3(N__13769),
            .lcout(\Lab_UT.scdp.key2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22622),
            .ce(),
            .sr(N__18056));
    defparam \Lab_UT.scdp.k3h.q_2_LC_7_14_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3h.q_2_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3h.q_2_LC_7_14_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.scdp.k3h.q_2_LC_7_14_2  (
            .in0(N__15559),
            .in1(N__15184),
            .in2(N__13815),
            .in3(N__13836),
            .lcout(\Lab_UT.scdp.key3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22622),
            .ce(),
            .sr(N__18056));
    defparam \Lab_UT.scdp.k3l.q_2_LC_7_14_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3l.q_2_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3l.q_2_LC_7_14_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k3l.q_2_LC_7_14_3  (
            .in0(N__15183),
            .in1(N__15560),
            .in2(N__13791),
            .in3(N__13724),
            .lcout(\Lab_UT.scdp.key3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22622),
            .ce(),
            .sr(N__18056));
    defparam \Lab_UT.scdp.k2h.q_3_LC_7_14_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2h.q_3_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2h.q_3_LC_7_14_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Lab_UT.scdp.k2h.q_3_LC_7_14_4  (
            .in0(N__13770),
            .in1(N__13740),
            .in2(N__15252),
            .in3(N__15323),
            .lcout(\Lab_UT.scdp.key2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22622),
            .ce(),
            .sr(N__18056));
    defparam \Lab_UT.scdp.k3l.q_3_LC_7_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3l.q_3_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3l.q_3_LC_7_14_5 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \Lab_UT.scdp.k3l.q_3_LC_7_14_5  (
            .in0(N__15321),
            .in1(N__13695),
            .in2(N__15248),
            .in3(N__13725),
            .lcout(\Lab_UT.scdp.key3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22622),
            .ce(),
            .sr(N__18056));
    defparam \Lab_UT.scctrl.state_ret_13_RNIHUNI41_LC_7_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNIHUNI41_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNIHUNI41_LC_7_14_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNIHUNI41_LC_7_14_6  (
            .in0(N__14194),
            .in1(N__14731),
            .in2(_gnd_net_),
            .in3(N__14980),
            .lcout(\Lab_UT.state_ret_13_RNIHUNI41_0 ),
            .ltout(\Lab_UT.state_ret_13_RNIHUNI41_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.k1l.q_2_LC_7_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1l.q_2_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1l.q_2_LC_7_14_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.scdp.k1l.q_2_LC_7_14_7  (
            .in0(N__15182),
            .in1(N__15557),
            .in2(N__14176),
            .in3(N__14169),
            .lcout(\Lab_UT.scdp.key1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22622),
            .ce(),
            .sr(N__18056));
    defparam \Lab_UT.scctrl.state_ret_8_RNIQ79K1_0_LC_7_15_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNIQ79K1_0_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNIQ79K1_0_LC_7_15_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNIQ79K1_0_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__14154),
            .in2(_gnd_net_),
            .in3(N__14119),
            .lcout(\Lab_UT.sccDnibble2En ),
            .ltout(\Lab_UT.sccDnibble2En_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_esr_RNO_2_LC_7_15_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_esr_RNO_2_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_esr_RNO_2_LC_7_15_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.scdp.u1.q_esr_RNO_2_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14104),
            .in3(N__14101),
            .lcout(\Lab_UT.scdp.u1.sccDnibble2En_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_1_LC_7_16_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_1_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u1.q_1_LC_7_16_6 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \Lab_UT.scdp.u1.q_1_LC_7_16_6  (
            .in0(N__14041),
            .in1(N__13988),
            .in2(_gnd_net_),
            .in3(N__14013),
            .lcout(\Lab_UT.scdp.byteToDecrypt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22616),
            .ce(),
            .sr(N__18060));
    defparam \Lab_UT.scctrl.next_state_2_LC_8_2_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_2_LC_8_2_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.next_state_2_LC_8_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scctrl.next_state_2_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13963),
            .lcout(\Lab_UT.scctrl.next_state_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22695),
            .ce(N__14792),
            .sr(N__18087));
    defparam \Lab_UT.scctrl.state_2_RNICEINI_2_LC_8_3_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNICEINI_2_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNICEINI_2_LC_8_3_0 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \Lab_UT.scctrl.state_2_RNICEINI_2_LC_8_3_0  (
            .in0(N__14218),
            .in1(N__18621),
            .in2(N__14233),
            .in3(N__18781),
            .lcout(\Lab_UT.scctrl.G_23_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIGC1Q_2_LC_8_3_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIGC1Q_2_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIGC1Q_2_LC_8_3_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIGC1Q_2_LC_8_3_1  (
            .in0(N__20081),
            .in1(N__19555),
            .in2(_gnd_net_),
            .in3(N__23065),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_i_a9_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_RNI7NLQ7_LC_8_3_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_RNI7NLQ7_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_11_RNI7NLQ7_LC_8_3_2 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_RNI7NLQ7_LC_8_3_2  (
            .in0(N__19163),
            .in1(N__20463),
            .in2(N__13918),
            .in3(N__22335),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_RNIK1DPL_LC_8_3_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_RNIK1DPL_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_11_RNIK1DPL_LC_8_3_3 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_RNIK1DPL_LC_8_3_3  (
            .in0(N__18623),
            .in1(N__14248),
            .in2(N__14242),
            .in3(N__14239),
            .lcout(\Lab_UT.scctrl.g0_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIU7GR_2_LC_8_3_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIU7GR_2_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIU7GR_2_LC_8_3_4 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIU7GR_2_LC_8_3_4  (
            .in0(N__19556),
            .in1(N__17497),
            .in2(N__20512),
            .in3(N__20079),
            .lcout(\Lab_UT.scctrl.G_23_0_a9_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_10_LC_8_3_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_10_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_10_LC_8_3_5 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_10_LC_8_3_5  (
            .in0(N__20080),
            .in1(N__22334),
            .in2(N__22065),
            .in3(N__20458),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_i_a10_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_8_LC_8_3_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_8_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_8_LC_8_3_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_8_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(N__18622),
            .in2(N__14221),
            .in3(N__18782),
            .lcout(\Lab_UT.scctrl.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNIGVQU8_LC_8_3_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNIGVQU8_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNIGVQU8_LC_8_3_7 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNIGVQU8_LC_8_3_7  (
            .in0(N__16003),
            .in1(N__20593),
            .in2(N__15997),
            .in3(N__19162),
            .lcout(\Lab_UT.scctrl.G_23_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNIK9N021_LC_8_4_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNIK9N021_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNIK9N021_LC_8_4_0 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNIK9N021_LC_8_4_0  (
            .in0(N__15914),
            .in1(N__15856),
            .in2(N__15897),
            .in3(N__15943),
            .lcout(\Lab_UT.scctrl.N_2ctr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIRRFK_LC_8_4_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIRRFK_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIRRFK_LC_8_4_1 .LUT_INIT=16'b0011001110110011;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNIRRFK_LC_8_4_1  (
            .in0(N__20091),
            .in1(N__17336),
            .in2(N__22422),
            .in3(N__21764),
            .lcout(\Lab_UT.scctrl.g0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_12_LC_8_4_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_12_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_12_LC_8_4_2 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_12_LC_8_4_2  (
            .in0(N__14302),
            .in1(N__14311),
            .in2(N__17095),
            .in3(N__14317),
            .lcout(\Lab_UT.state_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22685),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_9_LC_8_4_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_9_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_9_LC_8_4_3 .LUT_INIT=16'b0101011101011111;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_9_LC_8_4_3  (
            .in0(N__20089),
            .in1(N__21419),
            .in2(N__21172),
            .in3(N__21762),
            .lcout(\Lab_UT.scctrl.g0_i_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_LC_8_4_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_9_LC_8_4_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_LC_8_4_4  (
            .in0(N__14475),
            .in1(N__14347),
            .in2(_gnd_net_),
            .in3(N__14335),
            .lcout(\Lab_UT.un1_state_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22685),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIR10T_LC_8_4_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIR10T_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIR10T_LC_8_4_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep2_RNIR10T_LC_8_4_5  (
            .in0(N__20090),
            .in1(N__21420),
            .in2(N__22091),
            .in3(N__21763),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_23_0_a9_4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNIEA5S3_LC_8_4_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNIEA5S3_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNIEA5S3_LC_8_4_6 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNIEA5S3_LC_8_4_6  (
            .in0(N__21126),
            .in1(N__20092),
            .in2(N__14320),
            .in3(N__21023),
            .lcout(\Lab_UT.scctrl.G_23_0_3 ),
            .ltout(\Lab_UT.scctrl.G_23_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNIDDIN51_LC_8_4_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNIDDIN51_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNIDDIN51_LC_8_4_7 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNIDDIN51_LC_8_4_7  (
            .in0(N__14310),
            .in1(N__14301),
            .in2(N__14293),
            .in3(N__17091),
            .lcout(\Lab_UT.scctrl.N_3ctr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_16_LC_8_5_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_16_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_16_LC_8_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_16_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__20088),
            .in2(_gnd_net_),
            .in3(N__19237),
            .lcout(\Lab_UT.scctrl.g0_i_a7_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_RNILGT2_LC_8_5_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_RNILGT2_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_11_RNILGT2_LC_8_5_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_RNILGT2_LC_8_5_1  (
            .in0(_gnd_net_),
            .in1(N__22312),
            .in2(_gnd_net_),
            .in3(N__20443),
            .lcout(\Lab_UT.scctrl.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIGKQK_LC_8_5_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIGKQK_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIGKQK_LC_8_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNIGKQK_LC_8_5_2  (
            .in0(N__20442),
            .in1(N__22414),
            .in2(N__22333),
            .in3(N__23020),
            .lcout(\Lab_UT.scctrl.next_state_1_i_a5_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIS10T_LC_8_5_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIS10T_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIS10T_LC_8_5_3 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep1_RNIS10T_LC_8_5_3  (
            .in0(N__19293),
            .in1(N__21376),
            .in2(N__21128),
            .in3(N__21760),
            .lcout(\Lab_UT.scctrl.N_166_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_RNI7UQVB_LC_8_5_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNI7UQVB_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNI7UQVB_LC_8_5_4 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNI7UQVB_LC_8_5_4  (
            .in0(N__21869),
            .in1(N__14254),
            .in2(N__21202),
            .in3(N__20988),
            .lcout(\Lab_UT.scctrl.g0_0_i_2 ),
            .ltout(\Lab_UT.scctrl.g0_0_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_fast_LC_8_5_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_fast_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_8_fast_LC_8_5_5 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_fast_LC_8_5_5  (
            .in0(N__15896),
            .in1(N__15922),
            .in2(N__14446),
            .in3(N__15859),
            .lcout(\Lab_UT.scctrl.state_i_3_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22680),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_6_LC_8_5_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_6_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_6_LC_8_5_6 .LUT_INIT=16'b0011001000100000;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_6_LC_8_5_6  (
            .in0(N__21868),
            .in1(N__14410),
            .in2(N__21201),
            .in3(N__20987),
            .lcout(\Lab_UT.scctrl.g0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g1_1_o3_1_LC_8_5_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g1_1_o3_1_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g1_1_o3_1_LC_8_5_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Lab_UT.scdp.a2b.g1_1_o3_1_LC_8_5_7  (
            .in0(N__21377),
            .in1(N__21867),
            .in2(N__21129),
            .in3(N__21761),
            .lcout(\Lab_UT.scdp.a2b.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_0_RNI2GENA_1_LC_8_6_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_0_RNI2GENA_1_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_0_RNI2GENA_1_LC_8_6_0 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \Lab_UT.scctrl.state_0_RNI2GENA_1_LC_8_6_0  (
            .in0(N__21768),
            .in1(N__18599),
            .in2(N__16417),
            .in3(N__18772),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNI8MD1N_LC_8_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNI8MD1N_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNI8MD1N_LC_8_6_1 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNI8MD1N_LC_8_6_1  (
            .in0(N__14392),
            .in1(N__16009),
            .in2(N__14377),
            .in3(N__14374),
            .lcout(\Lab_UT.next_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep1_RNIP54M_LC_8_6_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep1_RNIP54M_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep1_RNIP54M_LC_8_6_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep1_RNIP54M_LC_8_6_2  (
            .in0(N__20062),
            .in1(N__19310),
            .in2(_gnd_net_),
            .in3(N__19238),
            .lcout(\Lab_UT.scctrl.G_21_i_a7_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIT10T_0_LC_8_6_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIT10T_0_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIT10T_0_LC_8_6_3 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep2_RNIT10T_0_LC_8_6_3  (
            .in0(N__21767),
            .in1(N__21161),
            .in2(N__22101),
            .in3(N__21401),
            .lcout(\Lab_UT.N_166_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI6J7KA_0_3_LC_8_6_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI6J7KA_0_3_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI6J7KA_0_3_LC_8_6_4 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI6J7KA_0_3_LC_8_6_4  (
            .in0(N__17482),
            .in1(N__19147),
            .in2(N__23064),
            .in3(N__20989),
            .lcout(\Lab_UT.scctrl.N_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_fast_LC_8_6_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_fast_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_13_fast_LC_8_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_fast_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20630),
            .lcout(\Lab_UT.scctrl.state_i_3_fast_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22675),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNI81K41_2_LC_8_6_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNI81K41_2_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNI81K41_2_LC_8_6_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNI81K41_2_LC_8_6_6  (
            .in0(N__19537),
            .in1(N__21765),
            .in2(_gnd_net_),
            .in3(N__22993),
            .lcout(\Lab_UT.scctrl.next_state_1_0_a5_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIT10T_LC_8_6_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIT10T_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIT10T_LC_8_6_7 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep2_RNIT10T_LC_8_6_7  (
            .in0(N__21766),
            .in1(N__21160),
            .in2(N__22100),
            .in3(N__21400),
            .lcout(\Lab_UT.scctrl.N_166_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.state_ret_5_rep2_RNIKU94_LC_8_7_0 .C_ON=1'b0;
    defparam \resetGen.state_ret_5_rep2_RNIKU94_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \resetGen.state_ret_5_rep2_RNIKU94_LC_8_7_0 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \resetGen.state_ret_5_rep2_RNIKU94_LC_8_7_0  (
            .in0(N__17616),
            .in1(N__18918),
            .in2(_gnd_net_),
            .in3(N__20051),
            .lcout(),
            .ltout(N_127_i_i_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNI2UI47_LC_8_7_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNI2UI47_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNI2UI47_LC_8_7_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNI2UI47_LC_8_7_1  (
            .in0(N__20930),
            .in1(N__21165),
            .in2(N__14509),
            .in3(N__14506),
            .lcout(\Lab_UT.scctrl.N_127_i_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_4_LC_8_7_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_4_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_4_LC_8_7_2 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_4_LC_8_7_2  (
            .in0(N__18355),
            .in1(N__16237),
            .in2(N__21195),
            .in3(N__20929),
            .lcout(\Lab_UT.scdp.a2b.g0_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g1_i_a4_0_2_LC_8_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g1_i_a4_0_2_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g1_i_a4_0_2_LC_8_7_3 .LUT_INIT=16'b1101000000000000;
    LogicCell40 \Lab_UT.scdp.a2b.g1_i_a4_0_2_LC_8_7_3  (
            .in0(N__20931),
            .in1(N__14497),
            .in2(N__17626),
            .in3(N__16669),
            .lcout(),
            .ltout(\Lab_UT.g1_i_a4_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNIRM5C62_LC_8_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNIRM5C62_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNIRM5C62_LC_8_7_4 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNIRM5C62_LC_8_7_4  (
            .in0(N__14491),
            .in1(N__16015),
            .in2(N__14485),
            .in3(N__16681),
            .lcout(),
            .ltout(\Lab_UT.g0_3_a3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_3_0_LC_8_7_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_3_0_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_3_0_LC_8_7_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Lab_UT.scdp.a2b.g0_3_0_LC_8_7_5  (
            .in0(N__14474),
            .in1(N__16378),
            .in2(N__14449),
            .in3(N__14551),
            .lcout(\Lab_UT.g0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIQB3N9_0_LC_8_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIQB3N9_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIQB3N9_0_LC_8_8_0 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIQB3N9_0_LC_8_8_0  (
            .in0(N__18749),
            .in1(N__14587),
            .in2(N__18600),
            .in3(N__23052),
            .lcout(\Lab_UT.N_182 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_12_LC_8_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_12_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_12_LC_8_8_1 .LUT_INIT=16'b0000101000101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_12_LC_8_8_1  (
            .in0(N__17494),
            .in1(N__18562),
            .in2(N__23089),
            .in3(N__18751),
            .lcout(\Lab_UT.scctrl.g0_1_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIQB3N9_0_0_LC_8_8_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIQB3N9_0_0_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIQB3N9_0_0_LC_8_8_2 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIQB3N9_0_0_LC_8_8_2  (
            .in0(N__18750),
            .in1(N__14566),
            .in2(N__18601),
            .in3(N__23053),
            .lcout(\Lab_UT.scctrl.N_182_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g1_i_a4_LC_8_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g1_i_a4_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g1_i_a4_LC_8_8_3 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \Lab_UT.scdp.a2b.g1_i_a4_LC_8_8_3  (
            .in0(N__21478),
            .in1(N__21529),
            .in2(N__17610),
            .in3(N__14537),
            .lcout(),
            .ltout(\Lab_UT.scdp.a2b.N_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_3_a3_0_3_LC_8_8_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_3_a3_0_3_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_3_a3_0_3_LC_8_8_4 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \Lab_UT.scdp.a2b.g0_3_a3_0_3_LC_8_8_4  (
            .in0(N__14713),
            .in1(N__14560),
            .in2(N__14554),
            .in3(N__17882),
            .lcout(\Lab_UT.scdp.a2b.g0_3_a3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIESKOU_3_LC_8_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIESKOU_3_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIESKOU_3_LC_8_8_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIESKOU_3_LC_8_8_5  (
            .in0(N__21477),
            .in1(N__21528),
            .in2(_gnd_net_),
            .in3(N__14536),
            .lcout(\Lab_UT.scctrl.next_state_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_a13_LC_8_8_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_a13_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_a13_LC_8_8_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_a13_LC_8_8_6  (
            .in0(N__19560),
            .in1(N__23051),
            .in2(N__16230),
            .in3(N__19090),
            .lcout(\Lab_UT.scdp.a2b.N_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIOBJ7V_3_LC_8_8_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIOBJ7V_3_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIOBJ7V_3_LC_8_8_7 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIOBJ7V_3_LC_8_8_7  (
            .in0(N__21479),
            .in1(N__21530),
            .in2(N__20282),
            .in3(N__14538),
            .lcout(\Lab_UT.scctrl.next_state_rst_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_3_LC_8_9_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_3_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_3_LC_8_9_0 .LUT_INIT=16'b1100101011111010;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_3_LC_8_9_0  (
            .in0(N__18325),
            .in1(N__16675),
            .in2(N__20093),
            .in3(N__14611),
            .lcout(\Lab_UT.scctrl.N_6_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNI3PVB9_2_LC_8_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNI3PVB9_2_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNI3PVB9_2_LC_8_9_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNI3PVB9_2_LC_8_9_1  (
            .in0(N__20530),
            .in1(N__18543),
            .in2(N__19553),
            .in3(N__18720),
            .lcout(\Lab_UT.state_2_RNI3PVB9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_14_LC_8_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_14_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_14_LC_8_9_2 .LUT_INIT=16'b1100110111111111;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_14_LC_8_9_2  (
            .in0(N__18719),
            .in1(N__19180),
            .in2(N__18589),
            .in3(N__21714),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_9_LC_8_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_9_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_9_LC_8_9_3 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_9_LC_8_9_3  (
            .in0(N__19679),
            .in1(_gnd_net_),
            .in2(N__14614),
            .in3(N__17476),
            .lcout(\Lab_UT.scctrl.g0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_3_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_3_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_3_LC_8_9_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_3_LC_8_9_4  (
            .in0(N__18982),
            .in1(N__14605),
            .in2(N__15013),
            .in3(N__14596),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_i_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_1_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_1_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_1_LC_8_9_5 .LUT_INIT=16'b0000010000001110;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_1_LC_8_9_5  (
            .in0(N__20052),
            .in1(N__20341),
            .in2(N__14590),
            .in3(N__18236),
            .lcout(\Lab_UT.scctrl.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNI1IP99_LC_8_9_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNI1IP99_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNI1IP99_LC_8_9_6 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNI1IP99_LC_8_9_6  (
            .in0(N__18721),
            .in1(N__19678),
            .in2(N__18590),
            .in3(N__21715),
            .lcout(\Lab_UT.scctrl.N_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI5GLD_3_LC_8_9_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI5GLD_3_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI5GLD_3_LC_8_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI5GLD_3_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__20487),
            .in2(_gnd_net_),
            .in3(N__17475),
            .lcout(\Lab_UT.scctrl.un6_sccDecrypt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNI67CB7_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNI67CB7_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNI67CB7_LC_8_10_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNI67CB7_LC_8_10_0  (
            .in0(N__21408),
            .in1(N__23062),
            .in2(_gnd_net_),
            .in3(N__19096),
            .lcout(\Lab_UT.scctrl.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIP9684_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIP9684_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIP9684_LC_8_10_1 .LUT_INIT=16'b1111111110001111;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep2_RNIP9684_LC_8_10_1  (
            .in0(N__22253),
            .in1(N__20537),
            .in2(N__22102),
            .in3(N__18729),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIRU4BD_LC_8_10_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIRU4BD_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIRU4BD_LC_8_10_2 .LUT_INIT=16'b1010100011111100;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep2_RNIRU4BD_LC_8_10_2  (
            .in0(N__16581),
            .in1(N__18572),
            .in2(N__14578),
            .in3(N__20990),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_RNIL9QO21_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNIL9QO21_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNIL9QO21_LC_8_10_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNIL9QO21_LC_8_10_3  (
            .in0(N__16693),
            .in1(N__14575),
            .in2(N__14569),
            .in3(N__17897),
            .lcout(\Lab_UT.scctrl.next_state_rst_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_RNIJN409_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_RNIJN409_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_11_RNIJN409_LC_8_10_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_RNIJN409_LC_8_10_4  (
            .in0(N__18728),
            .in1(N__20531),
            .in2(N__22304),
            .in3(N__18571),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_1_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIEANJ9_LC_8_10_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIEANJ9_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_RNIEANJ9_LC_8_10_5 .LUT_INIT=16'b0010001000101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep2_RNIEANJ9_LC_8_10_5  (
            .in0(N__17575),
            .in1(N__22096),
            .in2(N__14716),
            .in3(N__21189),
            .lcout(\Lab_UT.next_state_rst_1_3 ),
            .ltout(\Lab_UT.next_state_rst_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNO_0_0_LC_8_10_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNO_0_0_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNO_0_0_LC_8_10_6 .LUT_INIT=16'b0000111101001111;
    LogicCell40 \Lab_UT.scctrl.next_state_RNO_0_0_LC_8_10_6  (
            .in0(N__21409),
            .in1(N__23063),
            .in2(N__14704),
            .in3(N__19097),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_0_LC_8_10_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_0_LC_8_10_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.next_state_0_LC_8_10_7 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \Lab_UT.scctrl.next_state_0_LC_8_10_7  (
            .in0(N__20991),
            .in1(N__14700),
            .in2(N__14680),
            .in3(N__17898),
            .lcout(\Lab_UT.scctrl.next_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22648),
            .ce(N__14791),
            .sr(N__18084));
    defparam \Lab_UT.scctrl.state_ret_14_RNITPFM7_LC_8_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNITPFM7_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNITPFM7_LC_8_11_0 .LUT_INIT=16'b1111111100011111;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNITPFM7_LC_8_11_0  (
            .in0(N__23078),
            .in1(N__21397),
            .in2(N__21735),
            .in3(N__19101),
            .lcout(\Lab_UT.next_state_rst_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNIRVOO_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNIRVOO_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNIRVOO_LC_8_11_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNIRVOO_LC_8_11_1  (
            .in0(N__21398),
            .in1(N__21668),
            .in2(_gnd_net_),
            .in3(N__23079),
            .lcout(led_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_0_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_0_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_0_LC_8_11_2 .LUT_INIT=16'b0001000111110001;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_0_LC_8_11_2  (
            .in0(N__17218),
            .in1(N__14641),
            .in2(N__17119),
            .in3(N__17182),
            .lcout(\Lab_UT.scctrl.next_state_rst_0_3_N_6_1 ),
            .ltout(\Lab_UT.scctrl.next_state_rst_0_3_N_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_5_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_5_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_5_LC_8_11_3 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_5_LC_8_11_3  (
            .in0(N__20363),
            .in1(_gnd_net_),
            .in2(N__14629),
            .in3(N__14814),
            .lcout(\Lab_UT.scctrl.g0_i_m4_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_RNIOJNB3_LC_8_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNIOJNB3_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNIOJNB3_LC_8_11_4 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNIOJNB3_LC_8_11_4  (
            .in0(N__21196),
            .in1(N__21942),
            .in2(N__14752),
            .in3(N__21021),
            .lcout(\Lab_UT.scctrl.g0_i_2_0 ),
            .ltout(\Lab_UT.scctrl.g0_i_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_RNI3MOQ41_LC_8_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNI3MOQ41_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNI3MOQ41_LC_8_11_5 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNI3MOQ41_LC_8_11_5  (
            .in0(N__20364),
            .in1(N__14805),
            .in2(N__14626),
            .in3(N__17708),
            .lcout(\Lab_UT.scctrl.next_state_rst_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_1_LC_8_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_1_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.next_state_1_LC_8_11_6 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \Lab_UT.scctrl.next_state_1_LC_8_11_6  (
            .in0(N__17709),
            .in1(N__20365),
            .in2(N__14818),
            .in3(N__14806),
            .lcout(next_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22642),
            .ce(N__14794),
            .sr(N__18086));
    defparam \Lab_UT.scctrl.state_ret_14_RNI4BIC_LC_8_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNI4BIC_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNI4BIC_LC_8_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNI4BIC_LC_8_11_7  (
            .in0(N__21399),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21669),
            .lcout(\Lab_UT.scctrl.g0_i_a8_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep1_RNI2D76_LC_8_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep1_RNI2D76_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep1_RNI2D76_LC_8_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep1_RNI2D76_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__19834),
            .in2(_gnd_net_),
            .in3(N__19219),
            .lcout(\Lab_UT.scctrl.G_21_i_a7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_2_3_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_2_3_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_2_3_LC_8_12_1 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_2_3_LC_8_12_1  (
            .in0(N__17446),
            .in1(N__19107),
            .in2(N__23095),
            .in3(N__21022),
            .lcout(\Lab_UT.scctrl.N_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_1_3_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_1_3_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_1_3_LC_8_12_2 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_1_3_LC_8_12_2  (
            .in0(N__21688),
            .in1(N__18626),
            .in2(N__22801),
            .in3(N__18748),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_0_3_LC_8_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_0_3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_0_3_LC_8_12_3 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_0_3_LC_8_12_3  (
            .in0(N__19666),
            .in1(N__14743),
            .in2(N__14737),
            .in3(N__17442),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_1_0_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_3_LC_8_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_3_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_3_LC_8_12_4 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \Lab_UT.scctrl.state_1_3_LC_8_12_4  (
            .in0(N__18326),
            .in1(N__20284),
            .in2(N__14734),
            .in3(N__19835),
            .lcout(\Lab_UT.scctrl.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22636),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNI8TAR_LC_8_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNI8TAR_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNI8TAR_LC_8_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNI8TAR_LC_8_12_5  (
            .in0(N__20488),
            .in1(N__23086),
            .in2(N__19691),
            .in3(N__17441),
            .lcout(\Lab_UT.scctrl.next_state75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep1_LC_8_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep1_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_13_rep1_LC_8_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep1_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20631),
            .lcout(\Lab_UT.state_i_3_2_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22636),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_3_LC_8_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_3_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_3_LC_8_13_0 .LUT_INIT=16'b0000001010001010;
    LogicCell40 \Lab_UT.scctrl.state_ret_3_LC_8_13_0  (
            .in0(N__17731),
            .in1(N__19963),
            .in2(N__18332),
            .in3(N__17926),
            .lcout(\Lab_UT.scctrl.N_223_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22631),
            .ce(),
            .sr(N__18057));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_9_LC_8_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_9_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_9_LC_8_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_9_LC_8_13_1  (
            .in0(N__19961),
            .in1(N__18315),
            .in2(_gnd_net_),
            .in3(N__17367),
            .lcout(\Lab_UT.scctrl.N_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNO_3_LC_8_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_3_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_3_LC_8_13_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNO_3_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__18952),
            .in2(N__18331),
            .in3(N__19962),
            .lcout(\Lab_UT.scctrl.N_12_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_3_RNI95RN_LC_8_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_3_RNI95RN_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_3_RNI95RN_LC_8_13_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_3_RNI95RN_LC_8_13_3  (
            .in0(N__21769),
            .in1(N__23087),
            .in2(_gnd_net_),
            .in3(N__15001),
            .lcout(\Lab_UT.scctrl.next_state73 ),
            .ltout(\Lab_UT.scctrl.next_state73_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_3_RNII68F41_LC_8_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_3_RNII68F41_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_3_RNII68F41_LC_8_13_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \Lab_UT.scctrl.state_ret_3_RNII68F41_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__14908),
            .in2(N__14989),
            .in3(N__14981),
            .lcout(\Lab_UT.state_ret_3_RNII68F41_0 ),
            .ltout(\Lab_UT.state_ret_3_RNII68F41_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.k2l.q_0_LC_8_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2l.q_0_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2l.q_0_LC_8_13_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Lab_UT.scdp.k2l.q_0_LC_8_13_5  (
            .in0(N__15223),
            .in1(N__14943),
            .in2(N__14950),
            .in3(N__15511),
            .lcout(\Lab_UT.scdp.key2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22631),
            .ce(),
            .sr(N__18057));
    defparam \Lab_UT.scdp.k2l.q_1_LC_8_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2l.q_1_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2l.q_1_LC_8_13_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \Lab_UT.scdp.k2l.q_1_LC_8_13_6  (
            .in0(N__14928),
            .in1(N__15224),
            .in2(N__15390),
            .in3(N__14910),
            .lcout(\Lab_UT.scdp.key2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22631),
            .ce(),
            .sr(N__18057));
    defparam \Lab_UT.scdp.k2l.q_2_LC_8_13_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2l.q_2_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2l.q_2_LC_8_13_7 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Lab_UT.scdp.k2l.q_2_LC_8_13_7  (
            .in0(N__14909),
            .in1(N__14886),
            .in2(N__15273),
            .in3(N__15561),
            .lcout(\Lab_UT.scdp.key2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22631),
            .ce(),
            .sr(N__18057));
    defparam \Lab_UT.scdp.rxdataD.q_1_LC_8_14_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.rxdataD.q_1_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.rxdataD.q_1_LC_8_14_0 .LUT_INIT=16'b0100010111101111;
    LogicCell40 \Lab_UT.scdp.rxdataD.q_1_LC_8_14_0  (
            .in0(N__15819),
            .in1(N__15705),
            .in2(N__15789),
            .in3(N__14872),
            .lcout(\Lab_UT.scdp.binValD_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22627),
            .ce(),
            .sr(N__18059));
    defparam \Lab_UT.scdp.k0h.q_1_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0h.q_1_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0h.q_1_LC_8_14_1 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.scdp.k0h.q_1_LC_8_14_1  (
            .in0(N__15834),
            .in1(N__15364),
            .in2(N__15279),
            .in3(N__15430),
            .lcout(\Lab_UT.scdp.key0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22627),
            .ce(),
            .sr(N__18059));
    defparam \Lab_UT.scdp.rxdataD.q_2_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.rxdataD.q_2_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.rxdataD.q_2_LC_8_14_2 .LUT_INIT=16'b1111111101010000;
    LogicCell40 \Lab_UT.scdp.rxdataD.q_2_LC_8_14_2  (
            .in0(N__15820),
            .in1(_gnd_net_),
            .in2(N__15790),
            .in3(N__15706),
            .lcout(\Lab_UT.scdp.binValD_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22627),
            .ce(),
            .sr(N__18059));
    defparam \Lab_UT.scdp.k0h.q_2_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0h.q_2_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0h.q_2_LC_8_14_3 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \Lab_UT.scdp.k0h.q_2_LC_8_14_3  (
            .in0(N__15556),
            .in1(N__15528),
            .in2(N__15280),
            .in3(N__15431),
            .lcout(\Lab_UT.scdp.key0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22627),
            .ce(),
            .sr(N__18059));
    defparam \Lab_UT.scdp.k0h.q_0_LC_8_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0h.q_0_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0h.q_0_LC_8_14_5 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \Lab_UT.scdp.k0h.q_0_LC_8_14_5  (
            .in0(N__15510),
            .in1(N__15447),
            .in2(N__15278),
            .in3(N__15429),
            .lcout(\Lab_UT.scdp.key0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22627),
            .ce(),
            .sr(N__18059));
    defparam \Lab_UT.scdp.k0h.q_3_LC_8_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0h.q_3_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0h.q_3_LC_8_14_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k0h.q_3_LC_8_14_6  (
            .in0(N__15432),
            .in1(N__15324),
            .in2(N__15411),
            .in3(N__15265),
            .lcout(\Lab_UT.scdp.key0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22627),
            .ce(),
            .sr(N__18059));
    defparam \Lab_UT.scdp.k0l.q_1_LC_8_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0l.q_1_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0l.q_1_LC_8_14_7 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.scdp.k0l.q_1_LC_8_14_7  (
            .in0(N__15339),
            .in1(N__15365),
            .in2(N__15281),
            .in3(N__15077),
            .lcout(\Lab_UT.scdp.key0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22627),
            .ce(),
            .sr(N__18059));
    defparam \Lab_UT.scdp.k0l.q_3_LC_8_15_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0l.q_3_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0l.q_3_LC_8_15_7 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.scdp.k0l.q_3_LC_8_15_7  (
            .in0(N__15048),
            .in1(N__15325),
            .in2(N__15282),
            .in3(N__15082),
            .lcout(\Lab_UT.scdp.key0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22623),
            .ce(),
            .sr(N__18061));
    defparam \Lab_UT.scctrl.state_ret_13_RNIH6LF_LC_8_16_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNIH6LF_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNIH6LF_LC_8_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNIH6LF_LC_8_16_4  (
            .in0(N__21947),
            .in1(N__20538),
            .in2(N__19704),
            .in3(N__17498),
            .lcout(\Lab_UT.scctrl.next_state74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.state_ret_5_rep1_RNIP4DD_LC_9_3_1 .C_ON=1'b0;
    defparam \resetGen.state_ret_5_rep1_RNIP4DD_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \resetGen.state_ret_5_rep1_RNIP4DD_LC_9_3_1 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \resetGen.state_ret_5_rep1_RNIP4DD_LC_9_3_1  (
            .in0(N__20059),
            .in1(N__18938),
            .in2(N__17695),
            .in3(N__17359),
            .lcout(G_23_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIR2DQ_3_LC_9_3_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIR2DQ_3_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIR2DQ_3_LC_9_3_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIR2DQ_3_LC_9_3_5  (
            .in0(N__20454),
            .in1(N__23092),
            .in2(N__20094),
            .in3(N__17501),
            .lcout(\Lab_UT.scctrl.N_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNIOTIG_LC_9_4_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNIOTIG_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNIOTIG_LC_9_4_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNIOTIG_LC_9_4_0  (
            .in0(N__15984),
            .in1(N__19703),
            .in2(_gnd_net_),
            .in3(N__23093),
            .lcout(\Lab_UT.scctrl.g0_0_i_a8_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_RNI493D_LC_9_4_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNI493D_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNI493D_LC_9_4_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNI493D_LC_9_4_2  (
            .in0(N__21445),
            .in1(N__21870),
            .in2(_gnd_net_),
            .in3(N__21783),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_0_i_a8_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_RNIMMAAB_LC_9_4_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNIMMAAB_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNIMMAAB_LC_9_4_3 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNIMMAAB_LC_9_4_3  (
            .in0(N__15973),
            .in1(N__16024),
            .in2(N__15964),
            .in3(N__21024),
            .lcout(\Lab_UT.scctrl.g0_0_i_3_0 ),
            .ltout(\Lab_UT.scctrl.g0_0_i_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_LC_9_4_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_8_LC_9_4_4 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_LC_9_4_4  (
            .in0(N__15923),
            .in1(N__15891),
            .in2(N__15961),
            .in3(N__15944),
            .lcout(\Lab_UT.state_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22692),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_4_LC_9_4_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_4_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_4_LC_9_4_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_4_LC_9_4_5  (
            .in0(N__15958),
            .in1(N__16048),
            .in2(N__18954),
            .in3(N__15952),
            .lcout(\Lab_UT.scctrl.g0_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep2_LC_9_4_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_8_rep2_LC_9_4_6 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep2_LC_9_4_6  (
            .in0(N__15858),
            .in1(N__15895),
            .in2(N__15928),
            .in3(N__15946),
            .lcout(\Lab_UT.scctrl.state_i_3_0_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22692),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep1_LC_9_4_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_LC_9_4_7 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep1_LC_9_4_7  (
            .in0(N__15945),
            .in1(N__15924),
            .in2(N__15898),
            .in3(N__15857),
            .lcout(\Lab_UT.state_i_3_0_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22692),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNO_0_1_LC_9_5_0 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNO_0_1_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNO_0_1_LC_9_5_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ufifo.tx_fsm.cstate_RNO_0_1_LC_9_5_0  (
            .in0(N__20806),
            .in1(N__16207),
            .in2(N__16192),
            .in3(N__16170),
            .lcout(\ufifo.tx_fsm.N_60_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIR7JL_LC_9_5_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIR7JL_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIR7JL_LC_9_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep1_RNIR7JL_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__22378),
            .in2(_gnd_net_),
            .in3(N__19292),
            .lcout(\Lab_UT.scctrl.N_127_i_i_a6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_LC_9_5_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_LC_9_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20632),
            .lcout(\Lab_UT.state_i_3_2_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22686),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_7_LC_9_5_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_7_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_7_LC_9_5_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_7_LC_9_5_4  (
            .in0(N__19165),
            .in1(N__21388),
            .in2(N__23075),
            .in3(N__19970),
            .lcout(\Lab_UT.scctrl.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_RNIOI524_LC_9_5_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_RNIOI524_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_11_RNIOI524_LC_9_5_5 .LUT_INIT=16'b1010001000100010;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_RNIOI524_LC_9_5_5  (
            .in0(N__16042),
            .in1(N__22319),
            .in2(N__16036),
            .in3(N__20805),
            .lcout(\Lab_UT.scctrl.N_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNI73HE7_LC_9_5_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNI73HE7_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNI73HE7_LC_9_5_7 .LUT_INIT=16'b0101010101011101;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNI73HE7_LC_9_5_7  (
            .in0(N__17363),
            .in1(N__23022),
            .in2(N__21425),
            .in3(N__19164),
            .lcout(\Lab_UT.scctrl.g0_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIP81E9_LC_9_6_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIP81E9_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIP81E9_LC_9_6_0 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNIP81E9_LC_9_6_0  (
            .in0(N__21788),
            .in1(N__18624),
            .in2(N__22420),
            .in3(N__18783),
            .lcout(\Lab_UT.N_5 ),
            .ltout(\Lab_UT.N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_5_LC_9_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_5_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_5_LC_9_6_1 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_5_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__18367),
            .in2(N__16018),
            .in3(N__19161),
            .lcout(\Lab_UT.g0_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNIFT4T_LC_9_6_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNIFT4T_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNIFT4T_LC_9_6_3 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNIFT4T_LC_9_6_3  (
            .in0(N__20061),
            .in1(N__19697),
            .in2(N__17506),
            .in3(N__20229),
            .lcout(\Lab_UT.scctrl.g0_14_mb_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIDM3F1_LC_9_6_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIDM3F1_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIDM3F1_LC_9_6_5 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNIDM3F1_LC_9_6_5  (
            .in0(N__19538),
            .in1(N__22994),
            .in2(N__22069),
            .in3(N__22402),
            .lcout(\Lab_UT.scctrl.g0_0_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNI5UIN_LC_9_7_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNI5UIN_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNI5UIN_LC_9_7_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNI5UIN_LC_9_7_1  (
            .in0(N__20050),
            .in1(N__22407),
            .in2(N__22092),
            .in3(N__22259),
            .lcout(\Lab_UT.scctrl.N_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_8_LC_9_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_8_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_8_LC_9_7_3 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_8_LC_9_7_3  (
            .in0(N__19705),
            .in1(N__16393),
            .in2(N__16231),
            .in3(N__17524),
            .lcout(),
            .ltout(\Lab_UT.scdp.a2b.g0_iZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_3_LC_9_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_3_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_3_LC_9_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.scdp.a2b.g0_3_LC_9_7_4  (
            .in0(N__16387),
            .in1(N__16615),
            .in2(N__16381),
            .in3(N__16609),
            .lcout(\Lab_UT.scdp.a2b.g0_3_a3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.g0_i_a5_1_3_LC_9_7_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.g0_i_a5_1_3_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.g0_i_a5_1_3_LC_9_7_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.scctrl.g0_i_a5_1_3_LC_9_7_5  (
            .in0(N__16371),
            .in1(N__16970),
            .in2(N__16304),
            .in3(N__16560),
            .lcout(),
            .ltout(\Lab_UT.g0_i_a5_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_a13_2_LC_9_7_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_a13_2_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_a13_2_LC_9_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_a13_2_LC_9_7_6  (
            .in0(N__22406),
            .in1(N__19309),
            .in2(N__16240),
            .in3(N__20791),
            .lcout(\Lab_UT.scdp.a2b.N_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNO_7_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_7_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_7_LC_9_8_0 .LUT_INIT=16'b0101000100000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNO_7_LC_9_8_0  (
            .in0(N__20986),
            .in1(N__23011),
            .in2(N__19167),
            .in3(N__17490),
            .lcout(\Lab_UT.scctrl.N_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_o13_LC_9_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_o13_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_o13_LC_9_8_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_o13_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__22257),
            .in2(_gnd_net_),
            .in3(N__20539),
            .lcout(\Lab_UT.scdp.a2b.g1_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_4_LC_9_8_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_4_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_4_LC_9_8_2 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_4_LC_9_8_2  (
            .in0(N__16667),
            .in1(N__16213),
            .in2(N__20571),
            .in3(N__16603),
            .lcout(\Lab_UT.scctrl.g0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIPVJ8_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIPVJ8_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIPVJ8_LC_9_8_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNIPVJ8_LC_9_8_3  (
            .in0(N__22416),
            .in1(N__22258),
            .in2(_gnd_net_),
            .in3(N__20540),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_127_i_i_o6_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNI9IKA21_LC_9_8_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNI9IKA21_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNI9IKA21_LC_9_8_4 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNI9IKA21_LC_9_8_4  (
            .in0(N__17224),
            .in1(N__16624),
            .in2(N__16684),
            .in3(N__16605),
            .lcout(\Lab_UT.scctrl.N_127_i_i_a6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_8_LC_9_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_8_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_8_LC_9_8_5 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_8_LC_9_8_5  (
            .in0(N__17489),
            .in1(N__19151),
            .in2(N__23072),
            .in3(N__20985),
            .lcout(\Lab_UT.scctrl.N_190_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_9_LC_9_8_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_9_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_9_LC_9_8_6 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_9_LC_9_8_6  (
            .in0(N__16668),
            .in1(N__16642),
            .in2(N__16636),
            .in3(N__16623),
            .lcout(\Lab_UT.scdp.a2b.g0_iZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIDJ6UM_0_LC_9_8_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIDJ6UM_0_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIDJ6UM_0_LC_9_8_7 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIDJ6UM_0_LC_9_8_7  (
            .in0(N__16604),
            .in1(N__16588),
            .in2(N__16582),
            .in3(N__20984),
            .lcout(\Lab_UT.scctrl.g0_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNI0TTF2_LC_9_9_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNI0TTF2_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNI0TTF2_LC_9_9_0 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep1_RNI0TTF2_LC_9_9_0  (
            .in0(N__19314),
            .in1(N__16561),
            .in2(_gnd_net_),
            .in3(N__20758),
            .lcout(\Lab_UT.scctrl.next_state_1_i_o2_0_d_1 ),
            .ltout(\Lab_UT.scctrl.next_state_1_i_o2_0_d_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_1_LC_9_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_1_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_1_LC_9_9_1 .LUT_INIT=16'b0101000001110011;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_1_LC_9_9_1  (
            .in0(N__17170),
            .in1(N__17148),
            .in2(N__16513),
            .in3(N__17215),
            .lcout(\Lab_UT.state_ret_8_rep1_RNIJDTUE_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_rst_0_3_N_5L8_1_LC_9_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_rst_0_3_N_5L8_1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_rst_0_3_N_5L8_1_LC_9_9_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.scctrl.next_state_rst_0_3_N_5L8_1_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__16966),
            .in2(_gnd_net_),
            .in3(N__17076),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_0_3_N_5L8Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIKN433_LC_9_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIKN433_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIKN433_LC_9_9_3 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep1_RNIKN433_LC_9_9_3  (
            .in0(N__19315),
            .in1(N__16509),
            .in2(N__16450),
            .in3(N__16446),
            .lcout(\Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433 ),
            .ltout(\Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_LC_9_9_4 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_LC_9_9_4  (
            .in0(N__17149),
            .in1(N__17239),
            .in2(N__17227),
            .in3(N__17110),
            .lcout(\Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_7_LC_9_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_7_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_7_LC_9_9_5 .LUT_INIT=16'b0000101000111011;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_7_LC_9_9_5  (
            .in0(N__17111),
            .in1(N__17150),
            .in2(N__17178),
            .in3(N__17216),
            .lcout(\Lab_UT.scctrl.next_state_rst_0_3_N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_2_LC_9_9_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_2_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_2_LC_9_9_6 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_2_LC_9_9_6  (
            .in0(N__17217),
            .in1(N__17174),
            .in2(N__17155),
            .in3(N__17112),
            .lcout(\Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dk.shifter_ret_2_LC_9_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dk.shifter_ret_2_LC_9_9_7 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dk.shifter_ret_2_LC_9_9_7 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \Lab_UT.dk.shifter_ret_2_LC_9_9_7  (
            .in0(N__17077),
            .in1(_gnd_net_),
            .in2(N__16972),
            .in3(_gnd_net_),
            .lcout(resetGen_escKey_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22660),
            .ce(N__16759),
            .sr(N__18085));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_6_LC_9_10_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_6_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_6_LC_9_10_0 .LUT_INIT=16'b0100000011110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_6_LC_9_10_0  (
            .in0(N__21191),
            .in1(N__22435),
            .in2(N__17624),
            .in3(N__21015),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_2_LC_9_10_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_2_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_2_LC_9_10_1 .LUT_INIT=16'b1011000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_2_LC_9_10_1  (
            .in0(N__16729),
            .in1(N__16711),
            .in2(N__16705),
            .in3(N__16702),
            .lcout(\Lab_UT.scctrl.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIBABG4_2_LC_9_10_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIBABG4_2_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIBABG4_2_LC_9_10_2 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIBABG4_2_LC_9_10_2  (
            .in0(N__20569),
            .in1(N__17496),
            .in2(N__19554),
            .in3(N__18780),
            .lcout(\Lab_UT.scctrl.g0_i_a8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_8_RNI3O64_LC_9_10_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_8_RNI3O64_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_8_RNI3O64_LC_9_10_4 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \Lab_UT.scctrl.state_ret_8_RNI3O64_LC_9_10_4  (
            .in0(N__21190),
            .in1(N__17625),
            .in2(_gnd_net_),
            .in3(N__21922),
            .lcout(\Lab_UT.scctrl.g0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNITPFM7_0_LC_9_10_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNITPFM7_0_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNITPFM7_0_LC_9_10_5 .LUT_INIT=16'b1111111101010111;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNITPFM7_0_LC_9_10_5  (
            .in0(N__21756),
            .in1(N__23091),
            .in2(N__21444),
            .in3(N__19157),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_0_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNIB361N_LC_9_10_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNIB361N_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNIB361N_LC_9_10_6 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNIB361N_LC_9_10_6  (
            .in0(N__17611),
            .in1(N__17520),
            .in2(N__17509),
            .in3(N__18175),
            .lcout(\Lab_UT.scctrl.g0_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIT01T_3_LC_9_10_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIT01T_3_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIT01T_3_LC_9_10_7 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIT01T_3_LC_9_10_7  (
            .in0(N__17495),
            .in1(N__23090),
            .in2(N__17368),
            .in3(N__20570),
            .lcout(\Lab_UT.scctrl.g0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_2_LC_9_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_2_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_2_LC_9_11_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_2_LC_9_11_0  (
            .in0(N__18327),
            .in1(N__19877),
            .in2(_gnd_net_),
            .in3(N__18246),
            .lcout(\Lab_UT.scctrl.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNINBNBI_LC_9_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNINBNBI_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNINBNBI_LC_9_11_1 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNINBNBI_LC_9_11_1  (
            .in0(N__17752),
            .in1(N__17299),
            .in2(N__17293),
            .in3(N__18625),
            .lcout(\Lab_UT.scctrl.g0_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNITQ09E1_1_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNITQ09E1_1_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNITQ09E1_1_LC_9_11_2 .LUT_INIT=16'b0101111100110011;
    LogicCell40 \Lab_UT.scctrl.next_state_RNITQ09E1_1_LC_9_11_2  (
            .in0(N__17284),
            .in1(N__17681),
            .in2(N__17275),
            .in3(N__19876),
            .lcout(\Lab_UT.scctrl.g2 ),
            .ltout(\Lab_UT.scctrl.g2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIM7FBH2_0_LC_9_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIM7FBH2_0_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIM7FBH2_0_LC_9_11_3 .LUT_INIT=16'b0001000010110000;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIM7FBH2_0_LC_9_11_3  (
            .in0(N__19878),
            .in1(N__18422),
            .in2(N__17266),
            .in3(N__18102),
            .lcout(\Lab_UT.scctrl.N_223_1_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_0_LC_9_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_0_LC_9_11_4 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_0_LC_9_11_4  (
            .in0(N__19880),
            .in1(N__17263),
            .in2(N__17691),
            .in3(N__17257),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_222i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_LC_9_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_7_LC_9_11_5 .LUT_INIT=16'b1010101110101111;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_LC_9_11_5  (
            .in0(N__18922),
            .in1(N__17908),
            .in2(N__17248),
            .in3(N__17245),
            .lcout(Lab_UT_scctrl_N_221_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22649),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIDKJEO1_3_LC_9_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIDKJEO1_3_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIDKJEO1_3_LC_9_11_6 .LUT_INIT=16'b0000010010001100;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIDKJEO1_3_LC_9_11_6  (
            .in0(N__19879),
            .in1(N__17730),
            .in2(N__18336),
            .in3(N__17925),
            .lcout(\Lab_UT.scctrl.N_223_2_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_0_LC_9_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_0_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_0_LC_9_12_0 .LUT_INIT=16'b1111111100100111;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_0_LC_9_12_0  (
            .in0(N__19967),
            .in1(N__17902),
            .in2(N__18443),
            .in3(N__17863),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_i_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_LC_9_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_15_LC_9_12_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_LC_9_12_1  (
            .in0(N__17632),
            .in1(N__17851),
            .in2(N__17845),
            .in3(N__17716),
            .lcout(led_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22643),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNITPFM7_1_LC_9_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNITPFM7_1_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNITPFM7_1_LC_9_12_2 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNITPFM7_1_LC_9_12_2  (
            .in0(N__19149),
            .in1(N__21432),
            .in2(N__21792),
            .in3(N__23074),
            .lcout(\Lab_UT.scctrl.N_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIEUO38_2_LC_9_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIEUO38_2_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIEUO38_2_LC_9_12_3 .LUT_INIT=16'b0000010110001101;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIEUO38_2_LC_9_12_3  (
            .in0(N__19875),
            .in1(N__18346),
            .in2(N__20349),
            .in3(N__19148),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_18_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNIE2CTO_LC_9_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNIE2CTO_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNIE2CTO_LC_9_12_4 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNIE2CTO_LC_9_12_4  (
            .in0(N__19964),
            .in1(N__17743),
            .in2(N__17734),
            .in3(N__18802),
            .lcout(\Lab_UT.scctrl.next_stateZ0Z_2 ),
            .ltout(\Lab_UT.scctrl.next_stateZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_1_LC_9_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_1_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_1_LC_9_12_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_1_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__20267),
            .in2(N__17719),
            .in3(N__19966),
            .lcout(\Lab_UT.scctrl.N_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_15_RNO_3_LC_9_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_3_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_15_RNO_3_LC_9_12_6 .LUT_INIT=16'b1000110110101111;
    LogicCell40 \Lab_UT.scctrl.state_ret_15_RNO_3_LC_9_12_6  (
            .in0(N__19965),
            .in1(N__17710),
            .in2(N__17685),
            .in3(N__17638),
            .lcout(\Lab_UT.scctrl.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNI6VDS_0_2_LC_9_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNI6VDS_0_2_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNI6VDS_0_2_LC_9_13_0 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNI6VDS_0_2_LC_9_13_0  (
            .in0(N__19552),
            .in1(N__20574),
            .in2(N__22191),
            .in3(N__23077),
            .lcout(\Lab_UT.scctrl.g1_i_a7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_RNO_0_LC_9_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_RNO_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_11_RNO_0_LC_9_13_2 .LUT_INIT=16'b1100111101000111;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_RNO_0_LC_9_13_2  (
            .in0(N__20268),
            .in1(N__19968),
            .in2(N__18337),
            .in3(N__18247),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_LC_9_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_11_LC_9_13_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18223),
            .in3(N__18951),
            .lcout(\Lab_UT.state_i_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22637),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNI6VDS_2_LC_9_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNI6VDS_2_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNI6VDS_2_LC_9_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNI6VDS_2_LC_9_13_4  (
            .in0(N__19551),
            .in1(N__20572),
            .in2(N__22190),
            .in3(N__23076),
            .lcout(\Lab_UT.scctrl.next_state71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIR2DQ_2_LC_9_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIR2DQ_2_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIR2DQ_2_LC_9_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIR2DQ_2_LC_9_13_5  (
            .in0(N__19530),
            .in1(N__21943),
            .in2(N__22192),
            .in3(N__21770),
            .lcout(\Lab_UT.scctrl.next_state72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIPVJ8_0_LC_9_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIPVJ8_0_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIPVJ8_0_LC_9_13_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNIPVJ8_0_LC_9_13_6  (
            .in0(N__22415),
            .in1(N__22152),
            .in2(_gnd_net_),
            .in3(N__20573),
            .lcout(\Lab_UT.scctrl.g4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.EmsBitsSl_LC_9_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.EmsBitsSl_LC_9_14_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.EmsBitsSl_LC_9_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.scctrl.EmsBitsSl_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18140),
            .lcout(\Lab_UT.sccEmsBitsSl ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22632),
            .ce(),
            .sr(N__18062));
    defparam \Lab_UT.scctrl.state_ret_6_LC_9_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_6_LC_9_14_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_6_LC_9_14_7 .LUT_INIT=16'b0000001010001010;
    LogicCell40 \Lab_UT.scctrl.state_ret_6_LC_9_14_7  (
            .in0(N__18118),
            .in1(N__19969),
            .in2(N__18450),
            .in3(N__18109),
            .lcout(\Lab_UT.scctrl.N_223_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22632),
            .ce(),
            .sr(N__18062));
    defparam \Lab_UT.scctrl.state_1_RNO_5_0_LC_11_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_5_0_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_5_0_LC_11_6_1 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_5_0_LC_11_6_1  (
            .in0(N__21928),
            .in1(N__20565),
            .in2(N__22332),
            .in3(N__18784),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_0_i_a8_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_1_0_LC_11_6_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_1_0_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_1_0_LC_11_6_2 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_1_0_LC_11_6_2  (
            .in0(N__18379),
            .in1(N__18373),
            .in2(N__18472),
            .in3(N__18628),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_38_0_a3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_0_0_LC_11_6_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_0_0_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_0_0_LC_11_6_3 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_0_0_LC_11_6_3  (
            .in0(N__21562),
            .in1(N__18469),
            .in2(N__18454),
            .in3(N__21020),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_38_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_0_LC_11_6_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_0_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_0_LC_11_6_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Lab_UT.scctrl.state_1_0_LC_11_6_4  (
            .in0(N__18451),
            .in1(N__18869),
            .in2(N__18382),
            .in3(N__20070),
            .lcout(\Lab_UT.state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22687),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_6_0_LC_11_6_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_6_0_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_6_0_LC_11_6_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_6_0_LC_11_6_5  (
            .in0(N__21929),
            .in1(N__21185),
            .in2(_gnd_net_),
            .in3(N__21019),
            .lcout(\Lab_UT.scctrl.N_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_4_0_LC_11_6_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_4_0_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_4_0_LC_11_6_6 .LUT_INIT=16'b0000111100101111;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_4_0_LC_11_6_6  (
            .in0(N__22920),
            .in1(N__21407),
            .in2(N__20257),
            .in3(N__19156),
            .lcout(\Lab_UT.scctrl.g0_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_a9_1_0_LC_11_6_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_a9_1_0_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_a9_1_0_LC_11_6_7 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_a9_1_0_LC_11_6_7  (
            .in0(N__19521),
            .in1(N__20564),
            .in2(N__22331),
            .in3(N__22919),
            .lcout(\Lab_UT.scdp.a2b.g0_i_a9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_9_0_LC_11_7_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_9_0_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_9_0_LC_11_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_9_0_LC_11_7_0  (
            .in0(N__20556),
            .in1(N__19658),
            .in2(N__23019),
            .in3(N__22326),
            .lcout(\Lab_UT.scctrl.g0_0_i_a8_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_1_LC_11_7_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_1_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_1_LC_11_7_1 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_1_LC_11_7_1  (
            .in0(N__21975),
            .in1(N__18858),
            .in2(_gnd_net_),
            .in3(N__20019),
            .lcout(),
            .ltout(\Lab_UT.scdp.a2b.g0_iZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.g0_i_2_LC_11_7_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.g0_i_2_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.g0_i_2_LC_11_7_2 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \Lab_UT.scdp.a2b.g0_i_2_LC_11_7_2  (
            .in0(N__19319),
            .in1(N__22324),
            .in2(N__18358),
            .in3(N__19243),
            .lcout(\Lab_UT.scdp.a2b.g0_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_15_LC_11_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_15_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_15_LC_11_7_3 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_15_LC_11_7_3  (
            .in0(N__22323),
            .in1(N__20020),
            .in2(N__19323),
            .in3(N__20555),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_7_a13_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_12_LC_11_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_12_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_12_LC_11_7_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_12_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__18620),
            .in2(N__18973),
            .in3(N__18773),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_5_LC_11_7_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_5_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_5_LC_11_7_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_5_LC_11_7_5  (
            .in0(N__19371),
            .in1(N__19342),
            .in2(N__18970),
            .in3(N__18790),
            .lcout(\Lab_UT.scctrl.g0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_RNI7NLQ7_0_LC_11_7_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_RNI7NLQ7_0_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_11_RNI7NLQ7_0_LC_11_7_6 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_RNI7NLQ7_0_LC_11_7_6  (
            .in0(N__20554),
            .in1(N__22325),
            .in2(N__19393),
            .in3(N__19168),
            .lcout(\Lab_UT.scctrl.N_9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_0_LC_11_7_7 .C_ON=1'b0;
    defparam \resetGen.rst_0_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_0_LC_11_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_0_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22788),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22681),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIFKMJ3_LC_11_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIFKMJ3_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNIFKMJ3_LC_11_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNIFKMJ3_LC_11_8_0  (
            .in0(N__22421),
            .in1(N__18814),
            .in2(N__20815),
            .in3(N__22073),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_10_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNI0K8F7_LC_11_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNI0K8F7_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNI0K8F7_LC_11_8_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNI0K8F7_LC_11_8_1  (
            .in0(N__21961),
            .in1(N__21175),
            .in2(N__18805),
            .in3(N__20982),
            .lcout(\Lab_UT.scctrl.g1_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_13_LC_11_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_13_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_13_LC_11_8_3 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_13_LC_11_8_3  (
            .in0(N__19996),
            .in1(N__21174),
            .in2(N__22094),
            .in3(N__20981),
            .lcout(\Lab_UT.scctrl.N_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_0_RNIN6IE9_1_LC_11_8_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_0_RNIN6IE9_1_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_0_RNIN6IE9_1_LC_11_8_4 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \Lab_UT.scctrl.state_0_RNIN6IE9_1_LC_11_8_4  (
            .in0(N__21787),
            .in1(N__18765),
            .in2(N__18643),
            .in3(N__18616),
            .lcout(\Lab_UT.scctrl.N_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNIBRA17_LC_11_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNIBRA17_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNIBRA17_LC_11_8_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNIBRA17_LC_11_8_5  (
            .in0(N__19997),
            .in1(N__19429),
            .in2(N__21207),
            .in3(N__20983),
            .lcout(\Lab_UT.scctrl.G_21_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNO_0_LC_11_9_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_0_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_0_LC_11_9_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNO_0_LC_11_9_0  (
            .in0(N__19379),
            .in1(N__20270),
            .in2(_gnd_net_),
            .in3(N__19344),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_24_i_a4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_LC_11_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_14_LC_11_9_1 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_LC_11_9_1  (
            .in0(N__19408),
            .in1(N__21454),
            .in2(N__19396),
            .in3(N__20641),
            .lcout(\Lab_UT.N_169_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22667),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_2_LC_11_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_2_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_2_2_LC_11_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.scctrl.state_2_2_LC_11_9_2  (
            .in0(N__19381),
            .in1(N__19717),
            .in2(N__19360),
            .in3(N__19345),
            .lcout(\Lab_UT.state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22667),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIGC1Q_0_2_LC_11_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIGC1Q_0_2_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIGC1Q_0_2_LC_11_9_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIGC1Q_0_2_LC_11_9_3  (
            .in0(N__22955),
            .in1(N__19992),
            .in2(_gnd_net_),
            .in3(N__19486),
            .lcout(\Lab_UT.scctrl.G_21_i_a7_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNIPD53P_LC_11_9_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNIPD53P_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNIPD53P_LC_11_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNIPD53P_LC_11_9_4  (
            .in0(N__19380),
            .in1(N__19716),
            .in2(N__19359),
            .in3(N__19343),
            .lcout(\Lab_UT.scctrl.N_4ctr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_16_LC_11_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_16_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_16_LC_11_9_5 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_16_LC_11_9_5  (
            .in0(N__22956),
            .in1(N__19487),
            .in2(N__19327),
            .in3(N__19239),
            .lcout(\Lab_UT.scctrl.g0_1_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_15_LC_11_9_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_15_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_15_LC_11_9_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_15_LC_11_9_6  (
            .in0(N__19485),
            .in1(_gnd_net_),
            .in2(N__20069),
            .in3(N__22957),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_i_a7_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_10_LC_11_9_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_10_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_10_LC_11_9_7 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_10_LC_11_9_7  (
            .in0(N__22301),
            .in1(N__20578),
            .in2(N__19171),
            .in3(N__19155),
            .lcout(\Lab_UT.scctrl.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNO_4_LC_11_10_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_4_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_4_LC_11_10_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNO_4_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__21206),
            .in2(_gnd_net_),
            .in3(N__21025),
            .lcout(\Lab_UT.scctrl.N_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNO_8_LC_11_10_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_8_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_8_LC_11_10_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNO_8_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__19621),
            .in2(_gnd_net_),
            .in3(N__21948),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_24_i_o3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNO_5_LC_11_10_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_5_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_5_LC_11_10_3 .LUT_INIT=16'b1111100011111010;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNO_5_LC_11_10_3  (
            .in0(N__22297),
            .in1(N__20830),
            .in2(N__20818),
            .in3(N__20814),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_6_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNO_1_LC_11_10_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_1_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_1_LC_11_10_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNO_1_LC_11_10_4  (
            .in0(N__19972),
            .in1(N__20350),
            .in2(N__20650),
            .in3(N__20647),
            .lcout(\Lab_UT.scctrl.N_8_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_LC_11_10_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_13_LC_11_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20611),
            .lcout(\Lab_UT.state_i_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22663),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNIQT9P_LC_11_10_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNIQT9P_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNIQT9P_LC_11_10_6 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNIQT9P_LC_11_10_6  (
            .in0(N__19971),
            .in1(N__21290),
            .in2(N__21793),
            .in3(N__23002),
            .lcout(\Lab_UT.scctrl.G_23_0_a9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNI19C4_LC_11_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNI19C4_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNI19C4_LC_11_11_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNI19C4_LC_11_11_4  (
            .in0(N__22296),
            .in1(N__19628),
            .in2(_gnd_net_),
            .in3(N__20575),
            .lcout(\Lab_UT.scctrl.g0_i_a8_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIGKIO_2_LC_11_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIGKIO_2_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIGKIO_2_LC_11_11_5 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIGKIO_2_LC_11_11_5  (
            .in0(N__20348),
            .in1(N__20269),
            .in2(_gnd_net_),
            .in3(N__19998),
            .lcout(\Lab_UT.scctrl.G_21_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_3_3_LC_11_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_3_3_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_3_3_LC_11_12_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_3_3_LC_11_12_2  (
            .in0(N__19654),
            .in1(N__21951),
            .in2(N__19550),
            .in3(N__23018),
            .lcout(\Lab_UT.scctrl.g0_i_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.state_ret_5_fast_LC_12_7_2 .C_ON=1'b0;
    defparam \resetGen.state_ret_5_fast_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.state_ret_5_fast_LC_12_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \resetGen.state_ret_5_fast_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22789),
            .lcout(rst_i_3_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22688),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_7_RNO_13_LC_12_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_13_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_7_RNO_13_LC_12_7_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_7_RNO_13_LC_12_7_3  (
            .in0(N__21362),
            .in1(N__22077),
            .in2(_gnd_net_),
            .in3(N__21789),
            .lcout(\Lab_UT.scctrl.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNITKTS_LC_12_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNITKTS_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_rep2_RNITKTS_LC_12_7_4 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_rep2_RNITKTS_LC_12_7_4  (
            .in0(N__22423),
            .in1(N__22327),
            .in2(N__22095),
            .in3(N__21976),
            .lcout(\Lab_UT.scctrl.g1_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_3_0_LC_12_7_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_3_0_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_3_0_LC_12_7_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_3_0_LC_12_7_7  (
            .in0(N__21363),
            .in1(N__21923),
            .in2(N__21802),
            .in3(N__21790),
            .lcout(\Lab_UT.scctrl.state_1_RNO_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_14_RNO_2_LC_12_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_2_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_14_RNO_2_LC_12_8_5 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_14_RNO_2_LC_12_8_5  (
            .in0(N__21556),
            .in1(N__21547),
            .in2(N__21508),
            .in3(N__21490),
            .lcout(\Lab_UT.scctrl.N_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_6_RNIBMV1_LC_12_9_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_6_RNIBMV1_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_6_RNIBMV1_LC_12_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_6_RNIBMV1_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__21324),
            .in2(_gnd_net_),
            .in3(N__21253),
            .lcout(led_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // latticehx1k
