-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Jun 3 2019 04:43:08

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__23809\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \latticehx1k_pll_inst.clk\ : std_logic;
signal clk_in_c : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_1_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_0_cascade_\ : std_logic;
signal \buart.Z_tx.counter_RNIVE1P1_0_cascade_\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c3_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \ufifo_utb_txdata_rdy_0_i_1_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c2\ : std_logic;
signal ufifo_utb_txdata_rdy_0_i_1 : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.counter_RNIVE1P1_0\ : std_logic;
signal ufifo_fifo_txdata_6 : std_logic;
signal o_serial_data_c : std_logic;
signal \ufifo.fifo.fifo_txdata_7\ : std_logic;
signal \N_366_cascade_\ : std_logic;
signal \ufifo_utb_txdata_m0_7_cascade_\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal \ufifo.emitcrlf_fsm.cstate_ns_i_0_2_1_cascade_\ : std_logic;
signal \ufifo.N_323\ : std_logic;
signal \ufifo.emitcrlf_fsm.N_501_cascade_\ : std_logic;
signal \ufifo.emitcrlf_fsm.cstate_ns_i_0_0_1\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_0\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_1\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_2\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_3\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_4\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_5\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_6\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_7\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal ufifo_fifo_txdata_3 : std_logic;
signal \buart.Z_tx.N_369_cascade_\ : std_logic;
signal ufifo_fifo_txdata_4 : std_logic;
signal \buart.Z_tx.N_371_cascade_\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal \N_366\ : std_logic;
signal ufifo_fifo_txdata_5 : std_logic;
signal \buart.Z_tx.N_373_cascade_\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \buart.Z_tx.N_375\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal \buart.Z_tx.N_215_cascade_\ : std_logic;
signal \N_257_cascade_\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0_cascade_\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal \utb_txdata_1_cascade_\ : std_logic;
signal \N_257\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal \buart.Z_tx.N_58\ : std_logic;
signal ufifo_emitcrlf_fsm_cstate_0 : std_logic;
signal ufifo_emitcrlf_fsm_cstate_1 : std_logic;
signal \ufifo.fifo.wraddrZ0Z_2\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_3\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_7\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_8\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_0\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_1\ : std_logic;
signal \ufifo.tx_fsm.N_358_cascade_\ : std_logic;
signal \buart__tx_uart_busy_0\ : std_logic;
signal \ufifo.cstate_4\ : std_logic;
signal \ufifo.tx_fsm.N_394_cascade_\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_4\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_5\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_6\ : std_logic;
signal \ufifo.fifo.un1_emptyB_NE_0_cascade_\ : std_logic;
signal \ufifo.fifo.un1_emptyB_NE_3\ : std_logic;
signal \ufifo.fifo.un1_emptyB_NE_2\ : std_logic;
signal \ufifo.fifo.un1_emptyB_NE_4_cascade_\ : std_logic;
signal \ufifo.fifo.un1_emptyB_NE_1\ : std_logic;
signal \ufifo.emptyB_0_cascade_\ : std_logic;
signal \ufifo.tx_fsm.cstateZ0Z_5\ : std_logic;
signal \ufifo.tx_fsm.N_396_cascade_\ : std_logic;
signal \ufifo.tx_fsm.N_279\ : std_logic;
signal \ufifo.emptyB_0\ : std_logic;
signal \ufifo.tx_fsm.cstate_srsts_i_0_1_1_cascade_\ : std_logic;
signal \ufifo.tx_fsm.cstateZ0Z_1\ : std_logic;
signal \ufifo.fifo.fifo_txdata_2\ : std_logic;
signal \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0\ : std_logic;
signal \ufifo.sb_ram512x8_inst_RNILSN11_cascade_\ : std_logic;
signal utb_txdata_2 : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_rx.ser_clk\ : std_logic;
signal \buart.Z_rx.N_76_i\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_7\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_7\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_15\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.N_234_i_1_cascade_\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_23\ : std_logic;
signal \resetGen.N_421_cascade_\ : std_logic;
signal \buart.Z_tx.N_554\ : std_logic;
signal \resetGen.N_267_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \ufifo.popFifo\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_0\ : std_logic;
signal \bfn_4_4_0_\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_1\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_0\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_2\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_1\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_3\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_2\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_4\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_3\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_5\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_4\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_6\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_5\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_7\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_6\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_7\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_8\ : std_logic;
signal \N_251\ : std_logic;
signal \ufifo.fifo.fifo_txdata_1\ : std_logic;
signal \ufifo.sb_ram512x8_inst_RNIKRN11\ : std_logic;
signal ufifo_fifo_txdata_rdy : std_logic;
signal \buart.Z_tx.N_278\ : std_logic;
signal \resetGen.N_274\ : std_logic;
signal \resetGen.N_421\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal ufifo_tx_fsm_cstate_0 : std_logic;
signal \ufifo.fifo.fifo_txdata_0\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_0\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_1\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_2\ : std_logic;
signal \Lab_UT.scdp.b2a1.N_220_i_cascade_\ : std_logic;
signal \Lab_UT.scdp.b2a1.N_220_i\ : std_logic;
signal \Lab_UT.scdp.N_282_cascade_\ : std_logic;
signal \Lab_UT.scdp.b2a1.N_293\ : std_logic;
signal \Lab_UT.scctrl.sccLdLFSR\ : std_logic;
signal \Lab_UT.scctrl.EmsLoaded\ : std_logic;
signal \Lab_UT.scctrl.EmsLoaded_cascade_\ : std_logic;
signal \Lab_UT.sccElsBitsLd_cascade_\ : std_logic;
signal \Lab_UT.scdp.lsBits_i_1_6\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_6\ : std_logic;
signal \Lab_UT.scdp.N_282\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_6\ : std_logic;
signal \Lab_UT.scdp.b2a0.N_238_i_cascade_\ : std_logic;
signal \Lab_UT.scdp.b2a0.N_238_i\ : std_logic;
signal \Lab_UT.scdp.b2a0.N_227_i\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsD_6\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_5\ : std_logic;
signal \Lab_UT.scdp.b2a0.N_224_i\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsD_0\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_0\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsD_1\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_1\ : std_logic;
signal \Lab_UT.scdp.msBitsi.N_43_cascade_\ : std_logic;
signal \ufifo.txdataDZ0Z_1\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsD_2\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_2\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsD_4\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_4\ : std_logic;
signal \Lab_UT.scdp.lsBitsi.lsBitsDZ0Z_5\ : std_logic;
signal \Lab_UT.scdp.N_332_i_1_cascade_\ : std_logic;
signal \ufifo.txdataDZ0Z_5\ : std_logic;
signal \Lab_UT.sccEmsBitsSl\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsD_3\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_3\ : std_logic;
signal \Lab_UT.scdp.g0_0_i_1_0\ : std_logic;
signal \Lab_UT.scdp.msBitsi.N_1915_0\ : std_logic;
signal \ufifo.txdataDZ0Z_3\ : std_logic;
signal \Lab_UT.scdp.msBitsi.N_1919_0\ : std_logic;
signal \ufifo.txdataDZ0Z_2\ : std_logic;
signal \Lab_UT.scdp.msBitsi.N_1917_0\ : std_logic;
signal \ufifo.txdataDZ0Z_4\ : std_logic;
signal \Lab_UT.scdp.N_552\ : std_logic;
signal \Lab_UT.scdp.N_228_i_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.u0.byteToDecrypt_6\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.N_234_i_0\ : std_logic;
signal \Lab_UT.scdp.g0_0_i_1\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_0_1_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_225_i_0\ : std_logic;
signal \Lab_UT.scdp.u1.g0_0_i_a5_0_2_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_6\ : std_logic;
signal \Lab_UT.scdp.u1.g0_0_i_a5_0_2_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_6_0\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_0_a2_0_6\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_14\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30\ : std_logic;
signal \resetGen.N_243\ : std_logic;
signal \buart.bu_rx_data_i_2_4\ : std_logic;
signal \Lab_UT.scdp.msBitsi.q_esr_RNI679EZ0Z_6\ : std_logic;
signal \ufifo.txdataDZ0Z_6\ : std_logic;
signal \Lab_UT.scctrl.N_534\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_415_0\ : std_logic;
signal \Lab_UT.scctrl.g1_0_0\ : std_logic;
signal \Lab_UT.scctrl.g1_0_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_0_0_2_cascade_\ : std_logic;
signal \ufifo.txDataValidDZ0\ : std_logic;
signal \N_233_reti\ : std_logic;
signal \Lab_UT.scctrl.g1_0_1_0_cascade_\ : std_logic;
signal \Lab_UT.sccElsBitsLd\ : std_logic;
signal \Lab_UT.scdp.sccElsBitsLd_0\ : std_logic;
signal \Lab_UT.scctrl.g1_0_1_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_276\ : std_logic;
signal \Lab_UT.scdp.msBitsi.N_41\ : std_logic;
signal \ufifo.txdataDZ0Z_0\ : std_logic;
signal \Lab_UT.scctrl.N_46\ : std_logic;
signal \buart.Z_rx.sample_i_0_a2_0\ : std_logic;
signal \buart.Z_rx.N_230\ : std_logic;
signal \buart.Z_rx.N_230_cascade_\ : std_logic;
signal \Lab_UT.scdp.key0_7\ : std_logic;
signal \Lab_UT.scdp.key0_3\ : std_logic;
signal \Lab_UT.scdp.binVal_2_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_73\ : std_logic;
signal \Lab_UT.scdp.N_73_cascade_\ : std_logic;
signal \Lab_UT.scctrl.delayload\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_5_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_225_i_1\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21\ : std_logic;
signal \Lab_UT.scdp.u1.g0_0_i_a5_0_0_1_cascade_\ : std_logic;
signal \Lab_UT.scdp.u1.g0_0_i_a5_0_2_1\ : std_logic;
signal \Lab_UT.scdp.N_6_1\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_0_3_cascade_\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_3\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_3\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_0_3\ : std_logic;
signal \Lab_UT.scdp.N_226_i\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_0_1\ : std_logic;
signal \Lab_UT.scdp.u1.byteToDecrypt_1\ : std_logic;
signal \Lab_UT.scdp.u1.N_539_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_255_i\ : std_logic;
signal \Lab_UT.scdp.N_228_i\ : std_logic;
signal \Lab_UT.scdp.N_426_cascade_\ : std_logic;
signal \Lab_UT.scdp.q_RNI47LGA_1\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_4\ : std_logic;
signal \Lab_UT.scdp.b2a0.N_258_i\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_1_1\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_0_a2_0_4\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_0_a2_0_4_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_246_i\ : std_logic;
signal \Lab_UT.scdp.N_246_i_cascade_\ : std_logic;
signal \Lab_UT.scdp.u0.L4_tx_data_0_a2_1_6\ : std_logic;
signal \Lab_UT.scdp.N_256_i\ : std_logic;
signal \Lab_UT.scdp.key0_2\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_2_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_234_i\ : std_logic;
signal \Lab_UT.scdp.byteToDecrypt_5\ : std_logic;
signal \Lab_UT.scdp.N_228_i_0\ : std_logic;
signal \Lab_UT.scdp.g0_0_i_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_5\ : std_logic;
signal \Lab_UT.scdp.g0_0_i_1_1\ : std_logic;
signal \Lab_UT.scctrl.g1_1_1_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g2_0\ : std_logic;
signal \Lab_UT.scctrl.g1_3\ : std_logic;
signal \Lab_UT.scctrl.N_319_0\ : std_logic;
signal \Lab_UT.scctrl.N_414_0\ : std_logic;
signal \Lab_UT.scctrl.N_415_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1_0_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_259i\ : std_logic;
signal \Lab_UT.N_540i\ : std_logic;
signal \Lab_UT.scctrl.N_266\ : std_logic;
signal \Lab_UT.scctrl.N_472_0\ : std_logic;
signal \Lab_UT.scctrl.N_241_reti\ : std_logic;
signal \Lab_UT.scctrl.N_241_reti_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_263_0\ : std_logic;
signal \Lab_UT.scctrl.N_233_0\ : std_logic;
signal \Lab_UT.scctrl.N_351_1_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_5_1_cascade_\ : std_logic;
signal \CONSTANT_ONE_NET_cascade_\ : std_logic;
signal \ufifo.sb_ram512x8_inst_RNIKTQ21\ : std_logic;
signal \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1Z0Z_0\ : std_logic;
signal \N_368\ : std_logic;
signal utb_txdata_0 : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \buart.Z_rx.N_78\ : std_logic;
signal \Lab_UT.scctrl.N_418_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_2\ : std_logic;
signal \Lab_UT.scctrl.g0_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1_1\ : std_logic;
signal \Lab_UT.scctrl.N_418_2_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1_1_2\ : std_logic;
signal \Lab_UT.scctrl.N_39_i_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_22_i_cascade_\ : std_logic;
signal \Lab_UT.state_1_ret_0_RNI9C1NH_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.key3_5\ : std_logic;
signal \Lab_UT.state_1_ret_0_RNI9C1NH_0\ : std_logic;
signal \Lab_UT.scdp.key3_6\ : std_logic;
signal \Lab_UT.state_1_RNI6EDGH_0_2\ : std_logic;
signal \Lab_UT.scdp.key0_5\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_262_i\ : std_logic;
signal \Lab_UT.scdp.u1.g0_0_i_a5_0_0\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_0\ : std_logic;
signal \Lab_UT.scdp.u1.byteToDecryptZ0Z_2\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_2\ : std_logic;
signal \Lab_UT.scdp.u1.g0_0_i_a5_0_0_0\ : std_logic;
signal \Lab_UT.scdp.key0_6\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_6\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18\ : std_logic;
signal \Lab_UT.scdp.key0_4\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_4\ : std_logic;
signal \Lab_UT.scdp.key3_4\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_11\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_12\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9\ : std_logic;
signal \Lab_UT.sccLdLFSR_g\ : std_logic;
signal \Lab_UT.scctrl.N_534_reti_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_266i\ : std_logic;
signal bu_rx_data_2 : std_logic;
signal \Lab_UT.N_540\ : std_logic;
signal \Lab_UT.scctrl.N_399_0\ : std_logic;
signal \Lab_UT.scctrl.sccEldByte_i_a2_0Z0Z_1\ : std_logic;
signal \Lab_UT.scctrl.g2\ : std_logic;
signal \Lab_UT.scctrl.g1_0_5\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_0_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_444_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_319_1_0\ : std_logic;
signal \Lab_UT.scctrl.N_223_1_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_414_1_0\ : std_logic;
signal \Lab_UT.scctrl.N_444_0\ : std_logic;
signal \Lab_UT.scctrl.N_223_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_414_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1_0_2_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_0\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_1_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_5_1\ : std_logic;
signal \Lab_UT.scctrl.g0_2_0_0_a3_1_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_o7_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_12_2_cascade_\ : std_logic;
signal bu_rx_data_i_2_3_rep1 : std_logic;
signal \Lab_UT.scctrl.N_259\ : std_logic;
signal \Lab_UT.scctrl.g0_1_i_a8_0_1\ : std_logic;
signal \Lab_UT.scctrl.N_7_0\ : std_logic;
signal \Lab_UT.scctrl.N_10_0\ : std_logic;
signal \Lab_UT.scctrl.N_219\ : std_logic;
signal \buart__rx_shifter_0_fast_1\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0\ : std_logic;
signal \buart__rx_shifter_2_fast_6\ : std_logic;
signal \Lab_UT.scctrl.N_444\ : std_logic;
signal bu_rx_data_i_2_fast_3 : std_logic;
signal \N_243_reti\ : std_logic;
signal \Lab_UT.scctrl.N_219i\ : std_logic;
signal \Lab_UT.scctrl.N_271_0_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_1_cascade_\ : std_logic;
signal \buart__rx_shifter_0_fast_2\ : std_logic;
signal bu_rx_data_3 : std_logic;
signal \N_76_i_g\ : std_logic;
signal \buart.Z_rx.bitcountN11_15_i_0_o2_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_241\ : std_logic;
signal \Lab_UT.scctrl.g0_70_1_cascade_\ : std_logic;
signal \buart.Z_rx.N_80\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_2\ : std_logic;
signal \buart__rx_N_86_i_0_o2_1_0\ : std_logic;
signal \Lab_UT.N_252\ : std_logic;
signal \buart__rx_bitcount_4\ : std_logic;
signal \buart__rx_N_86_i_0_o2_1_0_cascade_\ : std_logic;
signal \buart__rx_bitcount_1\ : std_logic;
signal \Lab_UT.scctrl.r4.delay4\ : std_logic;
signal \Lab_UT.scctrl.delay3\ : std_logic;
signal \Lab_UT.scctrl.delay1\ : std_logic;
signal \Lab_UT.scctrl.delay2\ : std_logic;
signal \Lab_UT.scctrl.N_384\ : std_logic;
signal \Lab_UT.scctrl.N_385\ : std_logic;
signal \Lab_UT.scctrl.N_384_cascade_\ : std_logic;
signal \Lab_UT.N_100_i_cascade_\ : std_logic;
signal \Lab_UT.scdp.u2.N_100_i_0\ : std_logic;
signal \Lab_UT.scctrl.N_13_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_404_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_351\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_0_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_2\ : std_logic;
signal \Lab_UT.scctrl.N_6_2\ : std_logic;
signal \Lab_UT.scctrl.g0_8_1_0\ : std_logic;
signal \Lab_UT.scctrl.N_404_2\ : std_logic;
signal \Lab_UT.scctrl.g0_8_1_cascade_\ : std_logic;
signal \Lab_UT.scdp.key1_6\ : std_logic;
signal \Lab_UT.scdp.key1_7\ : std_logic;
signal \Lab_UT.scdp.key1_0\ : std_logic;
signal \Lab_UT.scdp.key1_3\ : std_logic;
signal \Lab_UT.scdp.key2_6\ : std_logic;
signal \Lab_UT.scdp.key2_4\ : std_logic;
signal \Lab_UT.scdp.key2_2\ : std_logic;
signal \Lab_UT.scdp.key1_2\ : std_logic;
signal \Lab_UT.scdp.key2_5\ : std_logic;
signal \Lab_UT.scdp.key1_4\ : std_logic;
signal \Lab_UT.scctrl.g1_0_4_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_3\ : std_logic;
signal \Lab_UT.scctrl.N_290_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_9_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_9_0\ : std_logic;
signal \Lab_UT.scctrl.g0_1_2_0\ : std_logic;
signal \Lab_UT.scctrl.g3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_1_4\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_i_0\ : std_logic;
signal \Lab_UT.scctrl.g3_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_7_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_10\ : std_logic;
signal \Lab_UT.scctrl.g0_1_i_0\ : std_logic;
signal \Lab_UT.scctrl.g0_1_i_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_1_i_4\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_2_0\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_a3_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_8\ : std_logic;
signal \Lab_UT.scctrl.N_290_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_8_3\ : std_logic;
signal \Lab_UT.scctrl.N_419_1\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_2_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_0_0\ : std_logic;
signal bu_rx_data_7 : std_logic;
signal \N_232\ : std_logic;
signal \Lab_UT.scctrl.g0_2_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_1_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_0_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_cascade_\ : std_logic;
signal \Lab_UT.scctrl.state_i_1_0_rep2\ : std_logic;
signal \Lab_UT.scctrl.N_299_i_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_4\ : std_logic;
signal \Lab_UT.scctrl.N_240_reti\ : std_logic;
signal \Lab_UT.scctrl.g0_2_0_0_a3_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_a3_3\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_a3_5_cascade_\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_a3_0_3\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_a3_0_1\ : std_logic;
signal \Lab_UT.scctrl.N_15\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_3_tz_0\ : std_logic;
signal \Lab_UT.scctrl.g0_0_4_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_4_1\ : std_logic;
signal \Lab_UT.scctrl.G_15_0_a10_1_2\ : std_logic;
signal \Lab_UT.scctrl.N_7\ : std_logic;
signal \Lab_UT.scctrl.g0_8_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_223_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_419_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_0_3\ : std_logic;
signal \Lab_UT.scctrl.N_418_1\ : std_logic;
signal \Lab_UT.scctrl.g0_8_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_8_2\ : std_logic;
signal \Lab_UT.scctrl.N_444_1\ : std_logic;
signal bu_rx_data_i_1_6 : std_logic;
signal bu_rx_data_4 : std_logic;
signal \Lab_UT.scctrl.G_24_i_a6_2_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_12_3\ : std_logic;
signal bu_rx_data_6 : std_logic;
signal \Lab_UT.scctrl.N_241_i_0\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_2_0\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_a6_0_2\ : std_logic;
signal \Lab_UT.scctrl.N_5_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_2_1\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_1_0\ : std_logic;
signal \Lab_UT.scctrl.N_401_0\ : std_logic;
signal \Lab_UT.scctrl.N_9_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_2\ : std_logic;
signal \Lab_UT.scctrl.N_170_i_cascade_\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_o6_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_17_i_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_20_i_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_277\ : std_logic;
signal \Lab_UT.scctrl.N_277_cascade_\ : std_logic;
signal \N_67\ : std_logic;
signal \Lab_UT.scctrl.N_355\ : std_logic;
signal \Lab_UT.scctrl.N_36\ : std_logic;
signal \Lab_UT.scctrl.N_27_i_cascade_\ : std_logic;
signal rst_i : std_logic;
signal \Lab_UT.scctrl.N_19\ : std_logic;
signal \Lab_UT.scctrl.N_415_2\ : std_logic;
signal \Lab_UT.scctrl.g1_2_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_stateZ0Z_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_2\ : std_logic;
signal \Lab_UT.scctrl.next_stateZ0Z_2\ : std_logic;
signal \Lab_UT.scctrl.g1_1_1_0\ : std_logic;
signal \Lab_UT.scctrl.g1_2_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_4_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_290_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_4_5\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_4_4_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_290_1\ : std_logic;
signal \Lab_UT.scctrl.g0_1_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_1_3\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_4_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_290\ : std_logic;
signal \Lab_UT.scctrl.next_state_0_3\ : std_logic;
signal \Lab_UT.scctrl.N_418_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1_0\ : std_logic;
signal \Lab_UT.scctrl.N_418\ : std_logic;
signal \Lab_UT.scctrl.N_415\ : std_logic;
signal \Lab_UT.scctrl.state_ret_0_fastZ0\ : std_logic;
signal \Lab_UT.scctrl.state_ret_4_RNOZ0Z_10_cascade_\ : std_logic;
signal \Lab_UT.scctrl.state_ret_4_RNOZ0Z_6\ : std_logic;
signal \Lab_UT.scctrl.N_295\ : std_logic;
signal \Lab_UT.scctrl.N_295_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_40_i\ : std_logic;
signal \Lab_UT.scctrl.N_487\ : std_logic;
signal \Lab_UT.scctrl.N_284\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_408_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a8_0_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_o7_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_12_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_408\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_3_tz\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_3_0_cascade_\ : std_logic;
signal rst_i_fast : std_logic;
signal \Lab_UT.scctrl.state_fast_3\ : std_logic;
signal \Lab_UT.scctrl.g0_0_0_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_0_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_0_3\ : std_logic;
signal \buart__rx_shifter_1_fast_0\ : std_logic;
signal \Lab_UT.scctrl.N_408_0\ : std_logic;
signal \Lab_UT.scctrl.g2_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_17\ : std_logic;
signal \Lab_UT.scctrl.N_240_i_0\ : std_logic;
signal bu_rx_data_i_1_5 : std_logic;
signal \Lab_UT.scctrl.N_412_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_1\ : std_logic;
signal \Lab_UT.scctrl.N_398i_i\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0_0\ : std_logic;
signal \Lab_UT.scctrl.nibbleInZ0Z1\ : std_logic;
signal \Lab_UT.scctrl.N_69_cascade_\ : std_logic;
signal \Lab_UT.sccDnibble1En_cascade_\ : std_logic;
signal \resetGen_rst_1_iso\ : std_logic;
signal \Lab_UT.scdp.u0.sccDnibble1En_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0dup_1\ : std_logic;
signal \Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93\ : std_logic;
signal \Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_69_i\ : std_logic;
signal \Lab_UT.scctrl.N_11\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst\ : std_logic;
signal \Lab_UT.scctrl.g0_9_a2_5_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1_1_0\ : std_logic;
signal \Lab_UT.scctrl.N_444_1_0\ : std_logic;
signal \Lab_UT.scctrl.g0_1_1\ : std_logic;
signal \Lab_UT.scctrl.g1_0_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1_2\ : std_logic;
signal \Lab_UT.scctrl.N_418_0_0\ : std_logic;
signal \Lab_UT.scctrl.g0_0\ : std_logic;
signal \Lab_UT.scctrl.g0_2_1\ : std_logic;
signal \Lab_UT.scctrl.g0_9_a2_2\ : std_logic;
signal \Lab_UT.scdp.byteToDecrypt_3\ : std_logic;
signal \Lab_UT.scdp.val_i_0_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.a2b.N_280\ : std_logic;
signal bu_rx_data_0 : std_logic;
signal \Lab_UT.scdp.N_378_cascade_\ : std_logic;
signal \Lab_UT.scdp.byteToDecrypt_4\ : std_logic;
signal \Lab_UT.scdp.val_i_0_0\ : std_logic;
signal \Lab_UT.scdp.N_378\ : std_logic;
signal \Lab_UT.scdp.u1.byteToDecryptZ0Z_0\ : std_logic;
signal \Lab_UT.scdp.a2b.val_0_tz_0_3\ : std_logic;
signal bu_rx_data_1 : std_logic;
signal bu_rx_data_i_2_2 : std_logic;
signal bu_rx_data_i_2_0 : std_logic;
signal \Lab_UT.sccDnibble1En\ : std_logic;
signal \Lab_UT.scdp.val_0_tz_3_cascade_\ : std_logic;
signal \Lab_UT.scdp.byteToDecrypt_7\ : std_logic;
signal \Lab_UT.scdp.key2_0\ : std_logic;
signal \Lab_UT.scdp.key2_1\ : std_logic;
signal \Lab_UT.scdp.key3_0\ : std_logic;
signal \Lab_UT.scdp.key3_1\ : std_logic;
signal \Lab_UT.scdp.binValD_2\ : std_logic;
signal \Lab_UT.scdp.key3_2\ : std_logic;
signal \Lab_UT.state_ret_12_RNIUVHQG_0\ : std_logic;
signal \Lab_UT.scdp.key3_3\ : std_logic;
signal \Lab_UT.scdp.val_0_tz_3\ : std_logic;
signal bu_rx_data_i_2_3 : std_logic;
signal \buart.Z_rx.N_301\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \buart__rx_hh_1\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \Lab_UT.scdp.binValD_0\ : std_logic;
signal \Lab_UT.scdp.key0_0\ : std_logic;
signal \Lab_UT.state_1_RNIO1RJH_0_2\ : std_logic;
signal \Lab_UT.scdp.key0_1\ : std_logic;
signal \Lab_UT.state_1_ret_3_RNI23U7H_0\ : std_logic;
signal \Lab_UT.scdp.key1_5\ : std_logic;
signal \Lab_UT.state_ret_RNIK5UKH_0\ : std_logic;
signal \Lab_UT.scdp.key2_3\ : std_logic;
signal \Lab_UT.scdp.binValD_1\ : std_logic;
signal \Lab_UT.state_ret_12_RNI2SEPG_0\ : std_logic;
signal \Lab_UT.scdp.key1_1\ : std_logic;
signal \Lab_UT.scdp.binVal_ValidD\ : std_logic;
signal \Lab_UT.scdp.binValD_3\ : std_logic;
signal \Lab_UT.state_1_RNI2IGHH_0_0\ : std_logic;
signal \Lab_UT.scdp.key2_7\ : std_logic;
signal \Lab_UT.scctrl.state_i_1_0\ : std_logic;
signal \Lab_UT.scctrl.N_296_i_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_RNO_1Z0Z_1\ : std_logic;
signal \Lab_UT.scctrl.N_319_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_1_0\ : std_logic;
signal \Lab_UT.scctrl.N_414_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_1_2\ : std_logic;
signal \Lab_UT.scctrl.N_319_1\ : std_logic;
signal \Lab_UT.scctrl.state_2_rep2\ : std_logic;
signal \Lab_UT.scctrl.N_7_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.G_18_i_a9_0_2\ : std_logic;
signal \Lab_UT.scctrl.G_18_i_1\ : std_logic;
signal \Lab_UT.scctrl.G_18_i_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.G_18_i_4_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_8_0_0\ : std_logic;
signal \Lab_UT.scctrl.g0_2_3_0\ : std_logic;
signal \Lab_UT.scctrl.g0_2_2_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_2_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_260_i_0\ : std_logic;
signal \Lab_UT.scctrl.N_404_4\ : std_logic;
signal bu_rx_data_5 : std_logic;
signal \Lab_UT.scctrl.g0_1_1_1\ : std_logic;
signal \Lab_UT.scctrl.g0_1_3\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_2_2\ : std_logic;
signal \Lab_UT.scctrl.N_13\ : std_logic;
signal \Lab_UT.scctrl.N_404_0\ : std_logic;
signal \Lab_UT.scctrl.N_5_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_12_0\ : std_logic;
signal \Lab_UT.scctrl.G_18_i_a9_0\ : std_logic;
signal \Lab_UT.scctrl.N_14_0\ : std_logic;
signal \Lab_UT.scctrl.stateZ0Z_2\ : std_logic;
signal \Lab_UT.scctrl.N_5\ : std_logic;
signal \Lab_UT.scctrl.N_21_0\ : std_logic;
signal \Lab_UT.scctrl.G_10_i_o7_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_a7_4_2\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_13_2\ : std_logic;
signal \Lab_UT.scctrl.rst_retZ0\ : std_logic;
signal \Lab_UT.scctrl.state_i_2_2\ : std_logic;
signal \Lab_UT.scctrl.N_12_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_8_0\ : std_logic;
signal \Lab_UT.scctrl.g0_9_a2_4\ : std_logic;
signal \Lab_UT.scctrl.state_3_rep1\ : std_logic;
signal \Lab_UT.scctrl.g0_9_a3_0_0\ : std_logic;
signal \Lab_UT.scctrl.next_stateZ0Z_3\ : std_logic;
signal \Lab_UT.scctrl.next_state_0_1\ : std_logic;
signal \Lab_UT.scctrl.m90_i_o6_0_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_404_1\ : std_logic;
signal \Lab_UT.scctrl.N_401\ : std_logic;
signal \Lab_UT.scctrl.N_399\ : std_logic;
signal \Lab_UT.scctrl.g0_2_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_2_3\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_356_1_0\ : std_logic;
signal \Lab_UT.scctrl.g0_9_a2_1\ : std_logic;
signal \Lab_UT.scctrl.g0_2_3_1\ : std_logic;
signal \Lab_UT.scctrl.next_stateZ0Z_0\ : std_logic;
signal \Lab_UT.scctrl.g0_2_2_1\ : std_logic;
signal rst : std_logic;
signal \Lab_UT.scctrl.next_state_3_0\ : std_logic;
signal \Lab_UT.scctrl.next_stateZ0Z_1\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_i_i_a2_1_0_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_6\ : std_logic;
signal \Lab_UT.scctrl.N_398\ : std_logic;
signal \Lab_UT.scctrl.N_235_i_0\ : std_logic;
signal \Lab_UT.scctrl.N_240\ : std_logic;
signal \Lab_UT.scctrl.N_296\ : std_logic;
signal \Lab_UT.scctrl.state_1_ret_1_RNICEVZ0Z81\ : std_logic;
signal \Lab_UT.scctrl.N_72_i_cascade_\ : std_logic;
signal \Lab_UT.state_ret_11_RNI4RQC3_0\ : std_logic;
signal \Lab_UT.state_ret_11_RNI4RQC3_0_cascade_\ : std_logic;
signal \N_74\ : std_logic;
signal \Lab_UT.sccDnibble2En\ : std_logic;
signal \Lab_UT.scctrl.N_223\ : std_logic;
signal \Lab_UT.scctrl.stateZ0Z_0\ : std_logic;
signal \Lab_UT.scctrl.N_5_0\ : std_logic;
signal \Lab_UT.scctrl.G_10_i_a7_0_2\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal clk_g : std_logic;
signal \Lab_UT.scctrl.next_state_RNIN96CP1Z0Z_3\ : std_logic;
signal \resetGen_rst_1_iso_g\ : std_logic;
signal \Lab_UT.scctrl.N_260\ : std_logic;
signal \Lab_UT.scctrl.N_235\ : std_logic;
signal \N_55_i\ : std_logic;
signal \Lab_UT.scctrl.state_i_1_0_rep1\ : std_logic;
signal \Lab_UT.scctrl.state_2_rep1\ : std_logic;
signal \Lab_UT.scctrl.N_13_1\ : std_logic;
signal \Lab_UT.scctrl.G_10_i_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.state_fast_2\ : std_logic;
signal \Lab_UT.scctrl.state_i_1_fast_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_0_2\ : std_logic;
signal rst_i_rep1 : std_logic;
signal \Lab_UT.scctrl.N_21_cascade_\ : std_logic;
signal \Lab_UT_scctrl_N_223_0\ : std_logic;
signal \N_272\ : std_logic;
signal \Lab_UT.scctrl.G_15_0_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.stateZ0Z_3\ : std_logic;
signal \Lab_UT.scctrl.G_15_0_2\ : std_logic;
signal \Lab_UT.scctrl.state_i_2_3\ : std_logic;
signal \N_21_1\ : std_logic;
signal \Lab_UT.scctrl.N_19_0\ : std_logic;
signal \Lab_UT.scctrl.N_8_1\ : std_logic;
signal \Lab_UT.scctrl.G_10_i_2\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_0_cascade_\ : std_logic;
signal rst_ii : std_logic;
signal \Lab_UT.scctrl.G_24_i_2\ : std_logic;
signal \Lab_UT.scctrl.N_273\ : std_logic;
signal \Lab_UT.scctrl.N_261\ : std_logic;
signal \Lab_UT.scctrl.stateZ0Z_1\ : std_logic;
signal \Lab_UT.scctrl.N_8_2\ : std_logic;
signal \Lab_UT.N_245\ : std_logic;
signal \N_245_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \ufifo.fifo.sb_ram512x8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \ufifo.fifo.sb_ram512x8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \ufifo.fifo.sb_ram512x8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \ufifo.fifo.sb_ram512x8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    led <= led_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    \ufifo.fifo.fifo_txdata_7\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(14);
    ufifo_fifo_txdata_6 <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(12);
    ufifo_fifo_txdata_5 <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(10);
    ufifo_fifo_txdata_4 <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(8);
    ufifo_fifo_txdata_3 <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(6);
    \ufifo.fifo.fifo_txdata_2\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(4);
    \ufifo.fifo.fifo_txdata_1\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(2);
    \ufifo.fifo.fifo_txdata_0\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(0);
    \ufifo.fifo.sb_ram512x8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__10293\&\N__10326\&\N__9897\&\N__9927\&\N__9957\&\N__9990\&\N__10023\&\N__10056\&\N__10086\;
    \ufifo.fifo.sb_ram512x8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__8979\&\N__9009\&\N__9399\&\N__9429\&\N__9456\&\N__9039\&\N__9066\&\N__8922\&\N__8949\;
    \ufifo.fifo.sb_ram512x8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \ufifo.fifo.sb_ram512x8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__11181\&'0'&\N__10848\&'0'&\N__10986\&'0'&\N__10758\&'0'&\N__11010\&'0'&\N__10914\&'0'&\N__11358\;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \ufifo.fifo.sb_ram512x8_inst_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\,
            RADDR => \ufifo.fifo.sb_ram512x8_inst_physical_RADDR_wire\,
            WADDR => \ufifo.fifo.sb_ram512x8_inst_physical_WADDR_wire\,
            MASK => \ufifo.fifo.sb_ram512x8_inst_physical_MASK_wire\,
            WDATA => \ufifo.fifo.sb_ram512x8_inst_physical_WDATA_wire\,
            RCLKE => \N__10140\,
            RCLK => \N__21135\,
            RE => \N__10130\,
            WCLKE => \N__11302\,
            WCLK => \N__21134\,
            WE => \N__11307\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \latticehx1k_pll_inst.clk\,
            REFERENCECLK => \N__8355\,
            RESETB => \N__21192\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23809\,
            DIN => \N__23808\,
            DOUT => \N__23807\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23809\,
            PADOUT => \N__23808\,
            PADIN => \N__23807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20541\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23800\,
            DIN => \N__23799\,
            DOUT => \N__23798\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23800\,
            PADOUT => \N__23799\,
            PADIN => \N__23798\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21588\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23791\,
            DIN => \N__23790\,
            DOUT => \N__23789\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23791\,
            PADOUT => \N__23790\,
            PADIN => \N__23789\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23782\,
            DIN => \N__23781\,
            DOUT => \N__23780\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23782\,
            PADOUT => \N__23781\,
            PADIN => \N__23780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21633\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23773\,
            DIN => \N__23772\,
            DOUT => \N__23771\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23773\,
            PADOUT => \N__23772\,
            PADIN => \N__23771\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__21114\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23764\,
            DIN => \N__23763\,
            DOUT => \N__23762\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__23764\,
            PADOUT => \N__23763\,
            PADIN => \N__23762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23755\,
            DIN => \N__23754\,
            DOUT => \N__23753\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23755\,
            PADOUT => \N__23754\,
            PADIN => \N__23753\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23746\,
            DIN => \N__23745\,
            DOUT => \N__23744\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23746\,
            PADOUT => \N__23745\,
            PADIN => \N__23744\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8562\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23737\,
            DIN => \N__23736\,
            DOUT => \N__23735\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23737\,
            PADOUT => \N__23736\,
            PADIN => \N__23735\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23728\,
            DIN => \N__23727\,
            DOUT => \N__23726\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23728\,
            PADOUT => \N__23727\,
            PADIN => \N__23726\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15525\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5815\ : CascadeMux
    port map (
            O => \N__23709\,
            I => \N__23701\
        );

    \I__5814\ : CascadeMux
    port map (
            O => \N__23708\,
            I => \N__23698\
        );

    \I__5813\ : CascadeMux
    port map (
            O => \N__23707\,
            I => \N__23692\
        );

    \I__5812\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23687\
        );

    \I__5811\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23676\
        );

    \I__5810\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23676\
        );

    \I__5809\ : InMux
    port map (
            O => \N__23701\,
            I => \N__23676\
        );

    \I__5808\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23676\
        );

    \I__5807\ : InMux
    port map (
            O => \N__23697\,
            I => \N__23676\
        );

    \I__5806\ : InMux
    port map (
            O => \N__23696\,
            I => \N__23673\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__23695\,
            I => \N__23669\
        );

    \I__5804\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23663\
        );

    \I__5803\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23663\
        );

    \I__5802\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23660\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__23687\,
            I => \N__23655\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__23676\,
            I => \N__23655\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__23673\,
            I => \N__23652\
        );

    \I__5798\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23649\
        );

    \I__5797\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23646\
        );

    \I__5796\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23643\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__23663\,
            I => \N__23638\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__23660\,
            I => \N__23638\
        );

    \I__5793\ : Span4Mux_h
    port map (
            O => \N__23655\,
            I => \N__23635\
        );

    \I__5792\ : Span4Mux_h
    port map (
            O => \N__23652\,
            I => \N__23630\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__23649\,
            I => \N__23630\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__23646\,
            I => \N__23625\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__23643\,
            I => \N__23625\
        );

    \I__5788\ : Span12Mux_s10_h
    port map (
            O => \N__23638\,
            I => \N__23622\
        );

    \I__5787\ : Span4Mux_v
    port map (
            O => \N__23635\,
            I => \N__23619\
        );

    \I__5786\ : Span4Mux_v
    port map (
            O => \N__23630\,
            I => \N__23614\
        );

    \I__5785\ : Span4Mux_s1_h
    port map (
            O => \N__23625\,
            I => \N__23614\
        );

    \I__5784\ : Odrv12
    port map (
            O => \N__23622\,
            I => \Lab_UT.scctrl.next_state_0_2\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__23619\,
            I => \Lab_UT.scctrl.next_state_0_2\
        );

    \I__5782\ : Odrv4
    port map (
            O => \N__23614\,
            I => \Lab_UT.scctrl.next_state_0_2\
        );

    \I__5781\ : InMux
    port map (
            O => \N__23607\,
            I => \N__23601\
        );

    \I__5780\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23596\
        );

    \I__5779\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23593\
        );

    \I__5778\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23590\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__23601\,
            I => \N__23586\
        );

    \I__5776\ : InMux
    port map (
            O => \N__23600\,
            I => \N__23581\
        );

    \I__5775\ : InMux
    port map (
            O => \N__23599\,
            I => \N__23581\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__23596\,
            I => \N__23574\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__23593\,
            I => \N__23574\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__23590\,
            I => \N__23574\
        );

    \I__5771\ : CascadeMux
    port map (
            O => \N__23589\,
            I => \N__23569\
        );

    \I__5770\ : Span4Mux_v
    port map (
            O => \N__23586\,
            I => \N__23564\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__23581\,
            I => \N__23564\
        );

    \I__5768\ : Span4Mux_s3_h
    port map (
            O => \N__23574\,
            I => \N__23561\
        );

    \I__5767\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23558\
        );

    \I__5766\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23553\
        );

    \I__5765\ : InMux
    port map (
            O => \N__23569\,
            I => \N__23553\
        );

    \I__5764\ : Span4Mux_v
    port map (
            O => \N__23564\,
            I => \N__23550\
        );

    \I__5763\ : Span4Mux_v
    port map (
            O => \N__23561\,
            I => \N__23547\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__23558\,
            I => \N__23544\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__23553\,
            I => \N__23535\
        );

    \I__5760\ : Span4Mux_s3_h
    port map (
            O => \N__23550\,
            I => \N__23535\
        );

    \I__5759\ : Span4Mux_s3_h
    port map (
            O => \N__23547\,
            I => \N__23535\
        );

    \I__5758\ : Span4Mux_v
    port map (
            O => \N__23544\,
            I => \N__23535\
        );

    \I__5757\ : Odrv4
    port map (
            O => \N__23535\,
            I => rst_i_rep1
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__23532\,
            I => \Lab_UT.scctrl.N_21_cascade_\
        );

    \I__5755\ : CascadeMux
    port map (
            O => \N__23529\,
            I => \N__23526\
        );

    \I__5754\ : InMux
    port map (
            O => \N__23526\,
            I => \N__23520\
        );

    \I__5753\ : InMux
    port map (
            O => \N__23525\,
            I => \N__23517\
        );

    \I__5752\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23514\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__23523\,
            I => \N__23510\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__23520\,
            I => \N__23484\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__23517\,
            I => \N__23481\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__23514\,
            I => \N__23478\
        );

    \I__5747\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23475\
        );

    \I__5746\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23470\
        );

    \I__5745\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23470\
        );

    \I__5744\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23467\
        );

    \I__5743\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23464\
        );

    \I__5742\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23458\
        );

    \I__5741\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23458\
        );

    \I__5740\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23455\
        );

    \I__5739\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23449\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__23502\,
            I => \N__23445\
        );

    \I__5737\ : CascadeMux
    port map (
            O => \N__23501\,
            I => \N__23435\
        );

    \I__5736\ : CascadeMux
    port map (
            O => \N__23500\,
            I => \N__23430\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__23499\,
            I => \N__23427\
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__23498\,
            I => \N__23422\
        );

    \I__5733\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23416\
        );

    \I__5732\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23416\
        );

    \I__5731\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23401\
        );

    \I__5730\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23401\
        );

    \I__5729\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23401\
        );

    \I__5728\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23401\
        );

    \I__5727\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23401\
        );

    \I__5726\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23401\
        );

    \I__5725\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23401\
        );

    \I__5724\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23398\
        );

    \I__5723\ : CascadeMux
    port map (
            O => \N__23487\,
            I => \N__23395\
        );

    \I__5722\ : Span4Mux_v
    port map (
            O => \N__23484\,
            I => \N__23381\
        );

    \I__5721\ : Span4Mux_v
    port map (
            O => \N__23481\,
            I => \N__23381\
        );

    \I__5720\ : Span4Mux_v
    port map (
            O => \N__23478\,
            I => \N__23381\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__23475\,
            I => \N__23378\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__23470\,
            I => \N__23373\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__23467\,
            I => \N__23373\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__23464\,
            I => \N__23370\
        );

    \I__5715\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23367\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__23458\,
            I => \N__23362\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__23455\,
            I => \N__23362\
        );

    \I__5712\ : InMux
    port map (
            O => \N__23454\,
            I => \N__23359\
        );

    \I__5711\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23356\
        );

    \I__5710\ : CascadeMux
    port map (
            O => \N__23452\,
            I => \N__23353\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__23449\,
            I => \N__23345\
        );

    \I__5708\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23334\
        );

    \I__5707\ : InMux
    port map (
            O => \N__23445\,
            I => \N__23334\
        );

    \I__5706\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23334\
        );

    \I__5705\ : InMux
    port map (
            O => \N__23443\,
            I => \N__23334\
        );

    \I__5704\ : InMux
    port map (
            O => \N__23442\,
            I => \N__23334\
        );

    \I__5703\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23323\
        );

    \I__5702\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23323\
        );

    \I__5701\ : InMux
    port map (
            O => \N__23439\,
            I => \N__23323\
        );

    \I__5700\ : InMux
    port map (
            O => \N__23438\,
            I => \N__23323\
        );

    \I__5699\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23323\
        );

    \I__5698\ : InMux
    port map (
            O => \N__23434\,
            I => \N__23318\
        );

    \I__5697\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23318\
        );

    \I__5696\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23305\
        );

    \I__5695\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23305\
        );

    \I__5694\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23305\
        );

    \I__5693\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23305\
        );

    \I__5692\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23305\
        );

    \I__5691\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23305\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__23416\,
            I => \N__23298\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__23401\,
            I => \N__23298\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__23398\,
            I => \N__23298\
        );

    \I__5687\ : InMux
    port map (
            O => \N__23395\,
            I => \N__23293\
        );

    \I__5686\ : InMux
    port map (
            O => \N__23394\,
            I => \N__23293\
        );

    \I__5685\ : InMux
    port map (
            O => \N__23393\,
            I => \N__23280\
        );

    \I__5684\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23280\
        );

    \I__5683\ : InMux
    port map (
            O => \N__23391\,
            I => \N__23280\
        );

    \I__5682\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23280\
        );

    \I__5681\ : InMux
    port map (
            O => \N__23389\,
            I => \N__23280\
        );

    \I__5680\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23280\
        );

    \I__5679\ : Span4Mux_v
    port map (
            O => \N__23381\,
            I => \N__23273\
        );

    \I__5678\ : Span4Mux_v
    port map (
            O => \N__23378\,
            I => \N__23273\
        );

    \I__5677\ : Span4Mux_v
    port map (
            O => \N__23373\,
            I => \N__23273\
        );

    \I__5676\ : Span4Mux_h
    port map (
            O => \N__23370\,
            I => \N__23264\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__23367\,
            I => \N__23264\
        );

    \I__5674\ : Span4Mux_s3_h
    port map (
            O => \N__23362\,
            I => \N__23264\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__23359\,
            I => \N__23264\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__23356\,
            I => \N__23261\
        );

    \I__5671\ : InMux
    port map (
            O => \N__23353\,
            I => \N__23252\
        );

    \I__5670\ : InMux
    port map (
            O => \N__23352\,
            I => \N__23252\
        );

    \I__5669\ : InMux
    port map (
            O => \N__23351\,
            I => \N__23252\
        );

    \I__5668\ : InMux
    port map (
            O => \N__23350\,
            I => \N__23252\
        );

    \I__5667\ : InMux
    port map (
            O => \N__23349\,
            I => \N__23247\
        );

    \I__5666\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23247\
        );

    \I__5665\ : Span4Mux_v
    port map (
            O => \N__23345\,
            I => \N__23242\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__23334\,
            I => \N__23242\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__23323\,
            I => \N__23239\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__23318\,
            I => \N__23230\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__23305\,
            I => \N__23230\
        );

    \I__5660\ : Span4Mux_v
    port map (
            O => \N__23298\,
            I => \N__23230\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__23293\,
            I => \N__23230\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__23280\,
            I => \Lab_UT_scctrl_N_223_0\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__23273\,
            I => \Lab_UT_scctrl_N_223_0\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__23264\,
            I => \Lab_UT_scctrl_N_223_0\
        );

    \I__5655\ : Odrv12
    port map (
            O => \N__23261\,
            I => \Lab_UT_scctrl_N_223_0\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__23252\,
            I => \Lab_UT_scctrl_N_223_0\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__23247\,
            I => \Lab_UT_scctrl_N_223_0\
        );

    \I__5652\ : Odrv4
    port map (
            O => \N__23242\,
            I => \Lab_UT_scctrl_N_223_0\
        );

    \I__5651\ : Odrv12
    port map (
            O => \N__23239\,
            I => \Lab_UT_scctrl_N_223_0\
        );

    \I__5650\ : Odrv4
    port map (
            O => \N__23230\,
            I => \Lab_UT_scctrl_N_223_0\
        );

    \I__5649\ : InMux
    port map (
            O => \N__23211\,
            I => \N__23203\
        );

    \I__5648\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23203\
        );

    \I__5647\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23199\
        );

    \I__5646\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23192\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__23203\,
            I => \N__23175\
        );

    \I__5644\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23172\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__23199\,
            I => \N__23169\
        );

    \I__5642\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23166\
        );

    \I__5641\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23163\
        );

    \I__5640\ : InMux
    port map (
            O => \N__23196\,
            I => \N__23157\
        );

    \I__5639\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23157\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__23192\,
            I => \N__23154\
        );

    \I__5637\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23151\
        );

    \I__5636\ : InMux
    port map (
            O => \N__23190\,
            I => \N__23144\
        );

    \I__5635\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23144\
        );

    \I__5634\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23141\
        );

    \I__5633\ : InMux
    port map (
            O => \N__23187\,
            I => \N__23138\
        );

    \I__5632\ : InMux
    port map (
            O => \N__23186\,
            I => \N__23129\
        );

    \I__5631\ : InMux
    port map (
            O => \N__23185\,
            I => \N__23129\
        );

    \I__5630\ : InMux
    port map (
            O => \N__23184\,
            I => \N__23129\
        );

    \I__5629\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23129\
        );

    \I__5628\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23123\
        );

    \I__5627\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23120\
        );

    \I__5626\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23112\
        );

    \I__5625\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23112\
        );

    \I__5624\ : InMux
    port map (
            O => \N__23178\,
            I => \N__23109\
        );

    \I__5623\ : Span4Mux_v
    port map (
            O => \N__23175\,
            I => \N__23105\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__23172\,
            I => \N__23100\
        );

    \I__5621\ : Span4Mux_v
    port map (
            O => \N__23169\,
            I => \N__23100\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__23166\,
            I => \N__23097\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__23163\,
            I => \N__23094\
        );

    \I__5618\ : InMux
    port map (
            O => \N__23162\,
            I => \N__23091\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__23157\,
            I => \N__23088\
        );

    \I__5616\ : Span4Mux_s3_h
    port map (
            O => \N__23154\,
            I => \N__23083\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__23151\,
            I => \N__23083\
        );

    \I__5614\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23080\
        );

    \I__5613\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23077\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__23144\,
            I => \N__23074\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__23141\,
            I => \N__23067\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__23138\,
            I => \N__23067\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__23129\,
            I => \N__23067\
        );

    \I__5608\ : InMux
    port map (
            O => \N__23128\,
            I => \N__23064\
        );

    \I__5607\ : InMux
    port map (
            O => \N__23127\,
            I => \N__23061\
        );

    \I__5606\ : InMux
    port map (
            O => \N__23126\,
            I => \N__23058\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__23123\,
            I => \N__23055\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__23120\,
            I => \N__23052\
        );

    \I__5603\ : InMux
    port map (
            O => \N__23119\,
            I => \N__23049\
        );

    \I__5602\ : InMux
    port map (
            O => \N__23118\,
            I => \N__23044\
        );

    \I__5601\ : InMux
    port map (
            O => \N__23117\,
            I => \N__23044\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__23112\,
            I => \N__23039\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__23109\,
            I => \N__23039\
        );

    \I__5598\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23036\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__23105\,
            I => \N__23023\
        );

    \I__5596\ : Span4Mux_v
    port map (
            O => \N__23100\,
            I => \N__23023\
        );

    \I__5595\ : Span4Mux_s2_h
    port map (
            O => \N__23097\,
            I => \N__23023\
        );

    \I__5594\ : Span4Mux_v
    port map (
            O => \N__23094\,
            I => \N__23023\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__23091\,
            I => \N__23023\
        );

    \I__5592\ : Span4Mux_v
    port map (
            O => \N__23088\,
            I => \N__23023\
        );

    \I__5591\ : Span4Mux_h
    port map (
            O => \N__23083\,
            I => \N__23010\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__23080\,
            I => \N__23010\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__23077\,
            I => \N__23010\
        );

    \I__5588\ : Span4Mux_v
    port map (
            O => \N__23074\,
            I => \N__23010\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__23067\,
            I => \N__23010\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__23064\,
            I => \N__23010\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__23061\,
            I => \N__23005\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__23058\,
            I => \N__23005\
        );

    \I__5583\ : Span4Mux_v
    port map (
            O => \N__23055\,
            I => \N__23000\
        );

    \I__5582\ : Span4Mux_s1_h
    port map (
            O => \N__23052\,
            I => \N__23000\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__23049\,
            I => \N__22993\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__23044\,
            I => \N__22993\
        );

    \I__5579\ : Span4Mux_h
    port map (
            O => \N__23039\,
            I => \N__22993\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__23036\,
            I => \N_272\
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__23023\,
            I => \N_272\
        );

    \I__5576\ : Odrv4
    port map (
            O => \N__23010\,
            I => \N_272\
        );

    \I__5575\ : Odrv4
    port map (
            O => \N__23005\,
            I => \N_272\
        );

    \I__5574\ : Odrv4
    port map (
            O => \N__23000\,
            I => \N_272\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__22993\,
            I => \N_272\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__22980\,
            I => \Lab_UT.scctrl.G_15_0_1_cascade_\
        );

    \I__5571\ : CascadeMux
    port map (
            O => \N__22977\,
            I => \N__22972\
        );

    \I__5570\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22958\
        );

    \I__5569\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22954\
        );

    \I__5568\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22951\
        );

    \I__5567\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22948\
        );

    \I__5566\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22945\
        );

    \I__5565\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22941\
        );

    \I__5564\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22934\
        );

    \I__5563\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22934\
        );

    \I__5562\ : InMux
    port map (
            O => \N__22966\,
            I => \N__22934\
        );

    \I__5561\ : InMux
    port map (
            O => \N__22965\,
            I => \N__22927\
        );

    \I__5560\ : InMux
    port map (
            O => \N__22964\,
            I => \N__22927\
        );

    \I__5559\ : InMux
    port map (
            O => \N__22963\,
            I => \N__22927\
        );

    \I__5558\ : InMux
    port map (
            O => \N__22962\,
            I => \N__22922\
        );

    \I__5557\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22922\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__22958\,
            I => \N__22919\
        );

    \I__5555\ : InMux
    port map (
            O => \N__22957\,
            I => \N__22915\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__22954\,
            I => \N__22912\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__22951\,
            I => \N__22909\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__22948\,
            I => \N__22906\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__22945\,
            I => \N__22903\
        );

    \I__5550\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22900\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__22941\,
            I => \N__22895\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__22934\,
            I => \N__22895\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__22927\,
            I => \N__22892\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__22922\,
            I => \N__22889\
        );

    \I__5545\ : Sp12to4
    port map (
            O => \N__22919\,
            I => \N__22885\
        );

    \I__5544\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22882\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__22915\,
            I => \N__22877\
        );

    \I__5542\ : Span4Mux_v
    port map (
            O => \N__22912\,
            I => \N__22877\
        );

    \I__5541\ : Span4Mux_v
    port map (
            O => \N__22909\,
            I => \N__22872\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__22906\,
            I => \N__22872\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__22903\,
            I => \N__22865\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__22900\,
            I => \N__22865\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__22895\,
            I => \N__22865\
        );

    \I__5536\ : Span4Mux_s2_h
    port map (
            O => \N__22892\,
            I => \N__22860\
        );

    \I__5535\ : Span4Mux_s2_h
    port map (
            O => \N__22889\,
            I => \N__22860\
        );

    \I__5534\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22857\
        );

    \I__5533\ : Odrv12
    port map (
            O => \N__22885\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__22882\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__22877\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__22872\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__5529\ : Odrv4
    port map (
            O => \N__22865\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__22860\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__22857\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__5526\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22836\
        );

    \I__5525\ : InMux
    port map (
            O => \N__22841\,
            I => \N__22836\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__22836\,
            I => \N__22833\
        );

    \I__5523\ : Odrv12
    port map (
            O => \N__22833\,
            I => \Lab_UT.scctrl.G_15_0_2\
        );

    \I__5522\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22816\
        );

    \I__5521\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22808\
        );

    \I__5520\ : InMux
    port map (
            O => \N__22828\,
            I => \N__22808\
        );

    \I__5519\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22808\
        );

    \I__5518\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22805\
        );

    \I__5517\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22793\
        );

    \I__5516\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22793\
        );

    \I__5515\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22793\
        );

    \I__5514\ : InMux
    port map (
            O => \N__22822\,
            I => \N__22793\
        );

    \I__5513\ : InMux
    port map (
            O => \N__22821\,
            I => \N__22785\
        );

    \I__5512\ : InMux
    port map (
            O => \N__22820\,
            I => \N__22782\
        );

    \I__5511\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22779\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__22816\,
            I => \N__22776\
        );

    \I__5509\ : InMux
    port map (
            O => \N__22815\,
            I => \N__22773\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__22808\,
            I => \N__22770\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__22805\,
            I => \N__22766\
        );

    \I__5506\ : InMux
    port map (
            O => \N__22804\,
            I => \N__22761\
        );

    \I__5505\ : InMux
    port map (
            O => \N__22803\,
            I => \N__22761\
        );

    \I__5504\ : InMux
    port map (
            O => \N__22802\,
            I => \N__22758\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__22793\,
            I => \N__22755\
        );

    \I__5502\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22752\
        );

    \I__5501\ : InMux
    port map (
            O => \N__22791\,
            I => \N__22747\
        );

    \I__5500\ : InMux
    port map (
            O => \N__22790\,
            I => \N__22747\
        );

    \I__5499\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22742\
        );

    \I__5498\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22742\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__22785\,
            I => \N__22738\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__22782\,
            I => \N__22733\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__22779\,
            I => \N__22730\
        );

    \I__5494\ : Span4Mux_s2_h
    port map (
            O => \N__22776\,
            I => \N__22723\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__22773\,
            I => \N__22723\
        );

    \I__5492\ : Span4Mux_h
    port map (
            O => \N__22770\,
            I => \N__22723\
        );

    \I__5491\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22720\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__22766\,
            I => \N__22717\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__22761\,
            I => \N__22714\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__22758\,
            I => \N__22707\
        );

    \I__5487\ : Span4Mux_s3_v
    port map (
            O => \N__22755\,
            I => \N__22707\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__22752\,
            I => \N__22707\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__22747\,
            I => \N__22704\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__22742\,
            I => \N__22701\
        );

    \I__5483\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22695\
        );

    \I__5482\ : Span4Mux_s2_h
    port map (
            O => \N__22738\,
            I => \N__22692\
        );

    \I__5481\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22687\
        );

    \I__5480\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22687\
        );

    \I__5479\ : Span12Mux_s6_h
    port map (
            O => \N__22733\,
            I => \N__22682\
        );

    \I__5478\ : Span12Mux_s10_v
    port map (
            O => \N__22730\,
            I => \N__22682\
        );

    \I__5477\ : Span4Mux_v
    port map (
            O => \N__22723\,
            I => \N__22679\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__22720\,
            I => \N__22670\
        );

    \I__5475\ : Span4Mux_s3_h
    port map (
            O => \N__22717\,
            I => \N__22670\
        );

    \I__5474\ : Span4Mux_v
    port map (
            O => \N__22714\,
            I => \N__22670\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__22707\,
            I => \N__22670\
        );

    \I__5472\ : Span4Mux_h
    port map (
            O => \N__22704\,
            I => \N__22665\
        );

    \I__5471\ : Span4Mux_s2_h
    port map (
            O => \N__22701\,
            I => \N__22665\
        );

    \I__5470\ : InMux
    port map (
            O => \N__22700\,
            I => \N__22658\
        );

    \I__5469\ : InMux
    port map (
            O => \N__22699\,
            I => \N__22658\
        );

    \I__5468\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22658\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__22695\,
            I => \Lab_UT.scctrl.state_i_2_3\
        );

    \I__5466\ : Odrv4
    port map (
            O => \N__22692\,
            I => \Lab_UT.scctrl.state_i_2_3\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__22687\,
            I => \Lab_UT.scctrl.state_i_2_3\
        );

    \I__5464\ : Odrv12
    port map (
            O => \N__22682\,
            I => \Lab_UT.scctrl.state_i_2_3\
        );

    \I__5463\ : Odrv4
    port map (
            O => \N__22679\,
            I => \Lab_UT.scctrl.state_i_2_3\
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__22670\,
            I => \Lab_UT.scctrl.state_i_2_3\
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__22665\,
            I => \Lab_UT.scctrl.state_i_2_3\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__22658\,
            I => \Lab_UT.scctrl.state_i_2_3\
        );

    \I__5459\ : InMux
    port map (
            O => \N__22641\,
            I => \N__22638\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__22638\,
            I => \N__22633\
        );

    \I__5457\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22630\
        );

    \I__5456\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22627\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__22633\,
            I => \N__22624\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__22630\,
            I => \N_21_1\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__22627\,
            I => \N_21_1\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__22624\,
            I => \N_21_1\
        );

    \I__5451\ : CascadeMux
    port map (
            O => \N__22617\,
            I => \N__22614\
        );

    \I__5450\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22611\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__22611\,
            I => \Lab_UT.scctrl.N_19_0\
        );

    \I__5448\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22605\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__22605\,
            I => \Lab_UT.scctrl.N_8_1\
        );

    \I__5446\ : InMux
    port map (
            O => \N__22602\,
            I => \N__22599\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__22599\,
            I => \Lab_UT.scctrl.G_10_i_2\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__22596\,
            I => \Lab_UT.scctrl.G_24_i_0_cascade_\
        );

    \I__5443\ : CascadeMux
    port map (
            O => \N__22593\,
            I => \N__22589\
        );

    \I__5442\ : CascadeMux
    port map (
            O => \N__22592\,
            I => \N__22586\
        );

    \I__5441\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22577\
        );

    \I__5440\ : InMux
    port map (
            O => \N__22586\,
            I => \N__22574\
        );

    \I__5439\ : InMux
    port map (
            O => \N__22585\,
            I => \N__22571\
        );

    \I__5438\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22564\
        );

    \I__5437\ : InMux
    port map (
            O => \N__22583\,
            I => \N__22564\
        );

    \I__5436\ : InMux
    port map (
            O => \N__22582\,
            I => \N__22564\
        );

    \I__5435\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22558\
        );

    \I__5434\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22555\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__22577\,
            I => \N__22552\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__22574\,
            I => \N__22549\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__22571\,
            I => \N__22543\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__22564\,
            I => \N__22543\
        );

    \I__5429\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22531\
        );

    \I__5428\ : InMux
    port map (
            O => \N__22562\,
            I => \N__22531\
        );

    \I__5427\ : InMux
    port map (
            O => \N__22561\,
            I => \N__22531\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__22558\,
            I => \N__22528\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__22555\,
            I => \N__22525\
        );

    \I__5424\ : Span4Mux_v
    port map (
            O => \N__22552\,
            I => \N__22520\
        );

    \I__5423\ : Span4Mux_s3_h
    port map (
            O => \N__22549\,
            I => \N__22520\
        );

    \I__5422\ : InMux
    port map (
            O => \N__22548\,
            I => \N__22517\
        );

    \I__5421\ : Span4Mux_s3_h
    port map (
            O => \N__22543\,
            I => \N__22514\
        );

    \I__5420\ : InMux
    port map (
            O => \N__22542\,
            I => \N__22511\
        );

    \I__5419\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22502\
        );

    \I__5418\ : InMux
    port map (
            O => \N__22540\,
            I => \N__22502\
        );

    \I__5417\ : InMux
    port map (
            O => \N__22539\,
            I => \N__22502\
        );

    \I__5416\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22502\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__22531\,
            I => \N__22499\
        );

    \I__5414\ : Span4Mux_h
    port map (
            O => \N__22528\,
            I => \N__22496\
        );

    \I__5413\ : Span4Mux_v
    port map (
            O => \N__22525\,
            I => \N__22493\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__22520\,
            I => \N__22490\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__22517\,
            I => \N__22485\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__22514\,
            I => \N__22485\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__22511\,
            I => rst_ii
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__22502\,
            I => rst_ii
        );

    \I__5407\ : Odrv12
    port map (
            O => \N__22499\,
            I => rst_ii
        );

    \I__5406\ : Odrv4
    port map (
            O => \N__22496\,
            I => rst_ii
        );

    \I__5405\ : Odrv4
    port map (
            O => \N__22493\,
            I => rst_ii
        );

    \I__5404\ : Odrv4
    port map (
            O => \N__22490\,
            I => rst_ii
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__22485\,
            I => rst_ii
        );

    \I__5402\ : InMux
    port map (
            O => \N__22470\,
            I => \N__22467\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__22467\,
            I => \Lab_UT.scctrl.G_24_i_2\
        );

    \I__5400\ : CascadeMux
    port map (
            O => \N__22464\,
            I => \N__22455\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__22463\,
            I => \N__22451\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__22462\,
            I => \N__22446\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__22461\,
            I => \N__22443\
        );

    \I__5396\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22437\
        );

    \I__5395\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22433\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__22458\,
            I => \N__22429\
        );

    \I__5393\ : InMux
    port map (
            O => \N__22455\,
            I => \N__22425\
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__22454\,
            I => \N__22421\
        );

    \I__5391\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22413\
        );

    \I__5390\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22413\
        );

    \I__5389\ : InMux
    port map (
            O => \N__22449\,
            I => \N__22413\
        );

    \I__5388\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22410\
        );

    \I__5387\ : InMux
    port map (
            O => \N__22443\,
            I => \N__22407\
        );

    \I__5386\ : InMux
    port map (
            O => \N__22442\,
            I => \N__22404\
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__22441\,
            I => \N__22401\
        );

    \I__5384\ : CascadeMux
    port map (
            O => \N__22440\,
            I => \N__22397\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__22437\,
            I => \N__22394\
        );

    \I__5382\ : InMux
    port map (
            O => \N__22436\,
            I => \N__22391\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__22433\,
            I => \N__22388\
        );

    \I__5380\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22383\
        );

    \I__5379\ : InMux
    port map (
            O => \N__22429\,
            I => \N__22383\
        );

    \I__5378\ : InMux
    port map (
            O => \N__22428\,
            I => \N__22380\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__22425\,
            I => \N__22377\
        );

    \I__5376\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22372\
        );

    \I__5375\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22372\
        );

    \I__5374\ : CascadeMux
    port map (
            O => \N__22420\,
            I => \N__22369\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__22413\,
            I => \N__22366\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__22410\,
            I => \N__22359\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__22407\,
            I => \N__22359\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__22404\,
            I => \N__22359\
        );

    \I__5369\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22356\
        );

    \I__5368\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22351\
        );

    \I__5367\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22351\
        );

    \I__5366\ : Span4Mux_h
    port map (
            O => \N__22394\,
            I => \N__22342\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__22391\,
            I => \N__22342\
        );

    \I__5364\ : Span4Mux_s1_h
    port map (
            O => \N__22388\,
            I => \N__22342\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__22383\,
            I => \N__22342\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__22380\,
            I => \N__22339\
        );

    \I__5361\ : Span4Mux_v
    port map (
            O => \N__22377\,
            I => \N__22334\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__22372\,
            I => \N__22334\
        );

    \I__5359\ : InMux
    port map (
            O => \N__22369\,
            I => \N__22331\
        );

    \I__5358\ : Span4Mux_h
    port map (
            O => \N__22366\,
            I => \N__22326\
        );

    \I__5357\ : Span4Mux_v
    port map (
            O => \N__22359\,
            I => \N__22326\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__22356\,
            I => \N__22323\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__22351\,
            I => \N__22316\
        );

    \I__5354\ : Span4Mux_v
    port map (
            O => \N__22342\,
            I => \N__22316\
        );

    \I__5353\ : Span4Mux_v
    port map (
            O => \N__22339\,
            I => \N__22316\
        );

    \I__5352\ : Sp12to4
    port map (
            O => \N__22334\,
            I => \N__22313\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__22331\,
            I => \N__22308\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__22326\,
            I => \N__22308\
        );

    \I__5349\ : Span4Mux_h
    port map (
            O => \N__22323\,
            I => \N__22303\
        );

    \I__5348\ : Span4Mux_h
    port map (
            O => \N__22316\,
            I => \N__22303\
        );

    \I__5347\ : Odrv12
    port map (
            O => \N__22313\,
            I => \Lab_UT.scctrl.N_273\
        );

    \I__5346\ : Odrv4
    port map (
            O => \N__22308\,
            I => \Lab_UT.scctrl.N_273\
        );

    \I__5345\ : Odrv4
    port map (
            O => \N__22303\,
            I => \Lab_UT.scctrl.N_273\
        );

    \I__5344\ : InMux
    port map (
            O => \N__22296\,
            I => \N__22293\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__22293\,
            I => \N__22281\
        );

    \I__5342\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22278\
        );

    \I__5341\ : InMux
    port map (
            O => \N__22291\,
            I => \N__22275\
        );

    \I__5340\ : InMux
    port map (
            O => \N__22290\,
            I => \N__22270\
        );

    \I__5339\ : InMux
    port map (
            O => \N__22289\,
            I => \N__22270\
        );

    \I__5338\ : InMux
    port map (
            O => \N__22288\,
            I => \N__22264\
        );

    \I__5337\ : InMux
    port map (
            O => \N__22287\,
            I => \N__22261\
        );

    \I__5336\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22251\
        );

    \I__5335\ : InMux
    port map (
            O => \N__22285\,
            I => \N__22251\
        );

    \I__5334\ : InMux
    port map (
            O => \N__22284\,
            I => \N__22247\
        );

    \I__5333\ : Span4Mux_v
    port map (
            O => \N__22281\,
            I => \N__22242\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__22278\,
            I => \N__22242\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__22275\,
            I => \N__22237\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22237\
        );

    \I__5329\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22230\
        );

    \I__5328\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22230\
        );

    \I__5327\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22227\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__22264\,
            I => \N__22224\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22221\
        );

    \I__5324\ : InMux
    port map (
            O => \N__22260\,
            I => \N__22210\
        );

    \I__5323\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22210\
        );

    \I__5322\ : InMux
    port map (
            O => \N__22258\,
            I => \N__22210\
        );

    \I__5321\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22210\
        );

    \I__5320\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22210\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__22251\,
            I => \N__22206\
        );

    \I__5318\ : InMux
    port map (
            O => \N__22250\,
            I => \N__22203\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__22247\,
            I => \N__22183\
        );

    \I__5316\ : Span4Mux_h
    port map (
            O => \N__22242\,
            I => \N__22178\
        );

    \I__5315\ : Span4Mux_s3_h
    port map (
            O => \N__22237\,
            I => \N__22178\
        );

    \I__5314\ : InMux
    port map (
            O => \N__22236\,
            I => \N__22170\
        );

    \I__5313\ : InMux
    port map (
            O => \N__22235\,
            I => \N__22170\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__22230\,
            I => \N__22165\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__22227\,
            I => \N__22165\
        );

    \I__5310\ : Span4Mux_v
    port map (
            O => \N__22224\,
            I => \N__22158\
        );

    \I__5309\ : Span4Mux_v
    port map (
            O => \N__22221\,
            I => \N__22158\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__22210\,
            I => \N__22158\
        );

    \I__5307\ : InMux
    port map (
            O => \N__22209\,
            I => \N__22155\
        );

    \I__5306\ : Span4Mux_h
    port map (
            O => \N__22206\,
            I => \N__22150\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__22203\,
            I => \N__22150\
        );

    \I__5304\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22141\
        );

    \I__5303\ : InMux
    port map (
            O => \N__22201\,
            I => \N__22141\
        );

    \I__5302\ : InMux
    port map (
            O => \N__22200\,
            I => \N__22141\
        );

    \I__5301\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22141\
        );

    \I__5300\ : InMux
    port map (
            O => \N__22198\,
            I => \N__22134\
        );

    \I__5299\ : InMux
    port map (
            O => \N__22197\,
            I => \N__22134\
        );

    \I__5298\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22134\
        );

    \I__5297\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22131\
        );

    \I__5296\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22126\
        );

    \I__5295\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22126\
        );

    \I__5294\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22123\
        );

    \I__5293\ : InMux
    port map (
            O => \N__22191\,
            I => \N__22116\
        );

    \I__5292\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22116\
        );

    \I__5291\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22116\
        );

    \I__5290\ : InMux
    port map (
            O => \N__22188\,
            I => \N__22109\
        );

    \I__5289\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22109\
        );

    \I__5288\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22109\
        );

    \I__5287\ : Span4Mux_v
    port map (
            O => \N__22183\,
            I => \N__22104\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__22178\,
            I => \N__22104\
        );

    \I__5285\ : InMux
    port map (
            O => \N__22177\,
            I => \N__22097\
        );

    \I__5284\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22097\
        );

    \I__5283\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22097\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__22170\,
            I => \N__22090\
        );

    \I__5281\ : Span4Mux_v
    port map (
            O => \N__22165\,
            I => \N__22090\
        );

    \I__5280\ : Span4Mux_h
    port map (
            O => \N__22158\,
            I => \N__22090\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__22155\,
            I => \N__22083\
        );

    \I__5278\ : Span4Mux_v
    port map (
            O => \N__22150\,
            I => \N__22083\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__22141\,
            I => \N__22083\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__22134\,
            I => \N__22076\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__22131\,
            I => \N__22076\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__22126\,
            I => \N__22076\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__22123\,
            I => \Lab_UT.scctrl.N_261\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__22116\,
            I => \Lab_UT.scctrl.N_261\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__22109\,
            I => \Lab_UT.scctrl.N_261\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__22104\,
            I => \Lab_UT.scctrl.N_261\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__22097\,
            I => \Lab_UT.scctrl.N_261\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__22090\,
            I => \Lab_UT.scctrl.N_261\
        );

    \I__5267\ : Odrv4
    port map (
            O => \N__22083\,
            I => \Lab_UT.scctrl.N_261\
        );

    \I__5266\ : Odrv12
    port map (
            O => \N__22076\,
            I => \Lab_UT.scctrl.N_261\
        );

    \I__5265\ : CascadeMux
    port map (
            O => \N__22059\,
            I => \N__22047\
        );

    \I__5264\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22038\
        );

    \I__5263\ : InMux
    port map (
            O => \N__22057\,
            I => \N__22024\
        );

    \I__5262\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22019\
        );

    \I__5261\ : InMux
    port map (
            O => \N__22055\,
            I => \N__22019\
        );

    \I__5260\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22016\
        );

    \I__5259\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22013\
        );

    \I__5258\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22010\
        );

    \I__5257\ : InMux
    port map (
            O => \N__22051\,
            I => \N__22003\
        );

    \I__5256\ : InMux
    port map (
            O => \N__22050\,
            I => \N__22003\
        );

    \I__5255\ : InMux
    port map (
            O => \N__22047\,
            I => \N__22003\
        );

    \I__5254\ : InMux
    port map (
            O => \N__22046\,
            I => \N__21998\
        );

    \I__5253\ : InMux
    port map (
            O => \N__22045\,
            I => \N__21998\
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__22044\,
            I => \N__21990\
        );

    \I__5251\ : InMux
    port map (
            O => \N__22043\,
            I => \N__21986\
        );

    \I__5250\ : InMux
    port map (
            O => \N__22042\,
            I => \N__21983\
        );

    \I__5249\ : InMux
    port map (
            O => \N__22041\,
            I => \N__21980\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__22038\,
            I => \N__21977\
        );

    \I__5247\ : InMux
    port map (
            O => \N__22037\,
            I => \N__21966\
        );

    \I__5246\ : InMux
    port map (
            O => \N__22036\,
            I => \N__21966\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__22035\,
            I => \N__21962\
        );

    \I__5244\ : InMux
    port map (
            O => \N__22034\,
            I => \N__21957\
        );

    \I__5243\ : InMux
    port map (
            O => \N__22033\,
            I => \N__21950\
        );

    \I__5242\ : InMux
    port map (
            O => \N__22032\,
            I => \N__21950\
        );

    \I__5241\ : InMux
    port map (
            O => \N__22031\,
            I => \N__21950\
        );

    \I__5240\ : CascadeMux
    port map (
            O => \N__22030\,
            I => \N__21945\
        );

    \I__5239\ : InMux
    port map (
            O => \N__22029\,
            I => \N__21938\
        );

    \I__5238\ : InMux
    port map (
            O => \N__22028\,
            I => \N__21938\
        );

    \I__5237\ : InMux
    port map (
            O => \N__22027\,
            I => \N__21938\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__22024\,
            I => \N__21929\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__21929\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__22016\,
            I => \N__21929\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__22013\,
            I => \N__21929\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__22010\,
            I => \N__21921\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__22003\,
            I => \N__21921\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__21998\,
            I => \N__21921\
        );

    \I__5229\ : InMux
    port map (
            O => \N__21997\,
            I => \N__21910\
        );

    \I__5228\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21910\
        );

    \I__5227\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21910\
        );

    \I__5226\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21910\
        );

    \I__5225\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21910\
        );

    \I__5224\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21905\
        );

    \I__5223\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21905\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__21986\,
            I => \N__21896\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__21983\,
            I => \N__21896\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21896\
        );

    \I__5219\ : Span4Mux_s2_v
    port map (
            O => \N__21977\,
            I => \N__21896\
        );

    \I__5218\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21889\
        );

    \I__5217\ : InMux
    port map (
            O => \N__21975\,
            I => \N__21889\
        );

    \I__5216\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21889\
        );

    \I__5215\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21882\
        );

    \I__5214\ : InMux
    port map (
            O => \N__21972\,
            I => \N__21882\
        );

    \I__5213\ : InMux
    port map (
            O => \N__21971\,
            I => \N__21882\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__21966\,
            I => \N__21879\
        );

    \I__5211\ : InMux
    port map (
            O => \N__21965\,
            I => \N__21876\
        );

    \I__5210\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21867\
        );

    \I__5209\ : InMux
    port map (
            O => \N__21961\,
            I => \N__21867\
        );

    \I__5208\ : InMux
    port map (
            O => \N__21960\,
            I => \N__21864\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__21957\,
            I => \N__21859\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__21950\,
            I => \N__21859\
        );

    \I__5205\ : CascadeMux
    port map (
            O => \N__21949\,
            I => \N__21855\
        );

    \I__5204\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21850\
        );

    \I__5203\ : InMux
    port map (
            O => \N__21945\,
            I => \N__21847\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__21938\,
            I => \N__21842\
        );

    \I__5201\ : Span4Mux_v
    port map (
            O => \N__21929\,
            I => \N__21842\
        );

    \I__5200\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21839\
        );

    \I__5199\ : Span4Mux_v
    port map (
            O => \N__21921\,
            I => \N__21836\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__21910\,
            I => \N__21831\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__21905\,
            I => \N__21831\
        );

    \I__5196\ : Span4Mux_v
    port map (
            O => \N__21896\,
            I => \N__21828\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__21889\,
            I => \N__21819\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__21882\,
            I => \N__21819\
        );

    \I__5193\ : Span4Mux_h
    port map (
            O => \N__21879\,
            I => \N__21819\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21819\
        );

    \I__5191\ : InMux
    port map (
            O => \N__21875\,
            I => \N__21809\
        );

    \I__5190\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21809\
        );

    \I__5189\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21809\
        );

    \I__5188\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21806\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__21867\,
            I => \N__21803\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__21864\,
            I => \N__21798\
        );

    \I__5185\ : Span4Mux_v
    port map (
            O => \N__21859\,
            I => \N__21798\
        );

    \I__5184\ : InMux
    port map (
            O => \N__21858\,
            I => \N__21795\
        );

    \I__5183\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21792\
        );

    \I__5182\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21787\
        );

    \I__5181\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21787\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__21850\,
            I => \N__21780\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21780\
        );

    \I__5178\ : Span4Mux_h
    port map (
            O => \N__21842\,
            I => \N__21780\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__21839\,
            I => \N__21775\
        );

    \I__5176\ : Span4Mux_h
    port map (
            O => \N__21836\,
            I => \N__21775\
        );

    \I__5175\ : Span4Mux_v
    port map (
            O => \N__21831\,
            I => \N__21768\
        );

    \I__5174\ : Span4Mux_h
    port map (
            O => \N__21828\,
            I => \N__21768\
        );

    \I__5173\ : Span4Mux_v
    port map (
            O => \N__21819\,
            I => \N__21768\
        );

    \I__5172\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21761\
        );

    \I__5171\ : InMux
    port map (
            O => \N__21817\,
            I => \N__21761\
        );

    \I__5170\ : InMux
    port map (
            O => \N__21816\,
            I => \N__21761\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__21809\,
            I => \N__21758\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__21806\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__21803\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__21798\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__21795\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__21792\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__21787\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5162\ : Odrv4
    port map (
            O => \N__21780\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5161\ : Odrv4
    port map (
            O => \N__21775\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__21768\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__21761\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5158\ : Odrv12
    port map (
            O => \N__21758\,
            I => \Lab_UT.scctrl.stateZ0Z_1\
        );

    \I__5157\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21732\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__21732\,
            I => \Lab_UT.scctrl.N_8_2\
        );

    \I__5155\ : CascadeMux
    port map (
            O => \N__21729\,
            I => \N__21725\
        );

    \I__5154\ : CascadeMux
    port map (
            O => \N__21728\,
            I => \N__21718\
        );

    \I__5153\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21714\
        );

    \I__5152\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21711\
        );

    \I__5151\ : CascadeMux
    port map (
            O => \N__21723\,
            I => \N__21703\
        );

    \I__5150\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21700\
        );

    \I__5149\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21697\
        );

    \I__5148\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21692\
        );

    \I__5147\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21692\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__21714\,
            I => \N__21687\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__21711\,
            I => \N__21687\
        );

    \I__5144\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21682\
        );

    \I__5143\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21682\
        );

    \I__5142\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21677\
        );

    \I__5141\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21677\
        );

    \I__5140\ : InMux
    port map (
            O => \N__21706\,
            I => \N__21672\
        );

    \I__5139\ : InMux
    port map (
            O => \N__21703\,
            I => \N__21672\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__21700\,
            I => \N__21669\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__21697\,
            I => \N__21666\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__21692\,
            I => \N__21663\
        );

    \I__5135\ : Span4Mux_v
    port map (
            O => \N__21687\,
            I => \N__21660\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__21682\,
            I => \N__21653\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__21677\,
            I => \N__21653\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__21672\,
            I => \N__21653\
        );

    \I__5131\ : Span4Mux_v
    port map (
            O => \N__21669\,
            I => \N__21650\
        );

    \I__5130\ : Span4Mux_h
    port map (
            O => \N__21666\,
            I => \N__21645\
        );

    \I__5129\ : Span4Mux_v
    port map (
            O => \N__21663\,
            I => \N__21645\
        );

    \I__5128\ : Sp12to4
    port map (
            O => \N__21660\,
            I => \N__21640\
        );

    \I__5127\ : Span12Mux_s8_v
    port map (
            O => \N__21653\,
            I => \N__21640\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__21650\,
            I => \Lab_UT.N_245\
        );

    \I__5125\ : Odrv4
    port map (
            O => \N__21645\,
            I => \Lab_UT.N_245\
        );

    \I__5124\ : Odrv12
    port map (
            O => \N__21640\,
            I => \Lab_UT.N_245\
        );

    \I__5123\ : IoInMux
    port map (
            O => \N__21633\,
            I => \N__21630\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__21630\,
            I => \N_245_i\
        );

    \I__5121\ : CascadeMux
    port map (
            O => \N__21627\,
            I => \Lab_UT.scctrl.N_72_i_cascade_\
        );

    \I__5120\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21615\
        );

    \I__5119\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21615\
        );

    \I__5118\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21615\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__21615\,
            I => \N__21612\
        );

    \I__5116\ : Span4Mux_v
    port map (
            O => \N__21612\,
            I => \N__21609\
        );

    \I__5115\ : Span4Mux_h
    port map (
            O => \N__21609\,
            I => \N__21605\
        );

    \I__5114\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21602\
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__21605\,
            I => \Lab_UT.state_ret_11_RNI4RQC3_0\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__21602\,
            I => \Lab_UT.state_ret_11_RNI4RQC3_0\
        );

    \I__5111\ : CascadeMux
    port map (
            O => \N__21597\,
            I => \Lab_UT.state_ret_11_RNI4RQC3_0_cascade_\
        );

    \I__5110\ : CascadeMux
    port map (
            O => \N__21594\,
            I => \N__21590\
        );

    \I__5109\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21585\
        );

    \I__5108\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21580\
        );

    \I__5107\ : InMux
    port map (
            O => \N__21589\,
            I => \N__21580\
        );

    \I__5106\ : IoInMux
    port map (
            O => \N__21588\,
            I => \N__21577\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__21585\,
            I => \N__21574\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__21580\,
            I => \N__21571\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__21577\,
            I => \N__21567\
        );

    \I__5102\ : Span4Mux_h
    port map (
            O => \N__21574\,
            I => \N__21562\
        );

    \I__5101\ : Span4Mux_h
    port map (
            O => \N__21571\,
            I => \N__21562\
        );

    \I__5100\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21558\
        );

    \I__5099\ : IoSpan4Mux
    port map (
            O => \N__21567\,
            I => \N__21555\
        );

    \I__5098\ : Span4Mux_h
    port map (
            O => \N__21562\,
            I => \N__21552\
        );

    \I__5097\ : InMux
    port map (
            O => \N__21561\,
            I => \N__21549\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__21558\,
            I => \N__21546\
        );

    \I__5095\ : Odrv4
    port map (
            O => \N__21555\,
            I => \N_74\
        );

    \I__5094\ : Odrv4
    port map (
            O => \N__21552\,
            I => \N_74\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__21549\,
            I => \N_74\
        );

    \I__5092\ : Odrv4
    port map (
            O => \N__21546\,
            I => \N_74\
        );

    \I__5091\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21531\
        );

    \I__5090\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21531\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__21531\,
            I => \N__21528\
        );

    \I__5088\ : Span4Mux_h
    port map (
            O => \N__21528\,
            I => \N__21525\
        );

    \I__5087\ : Odrv4
    port map (
            O => \N__21525\,
            I => \Lab_UT.sccDnibble2En\
        );

    \I__5086\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21515\
        );

    \I__5085\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21511\
        );

    \I__5084\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21508\
        );

    \I__5083\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21503\
        );

    \I__5082\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21503\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__21515\,
            I => \N__21492\
        );

    \I__5080\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21489\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__21511\,
            I => \N__21484\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__21508\,
            I => \N__21484\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__21503\,
            I => \N__21481\
        );

    \I__5076\ : InMux
    port map (
            O => \N__21502\,
            I => \N__21472\
        );

    \I__5075\ : InMux
    port map (
            O => \N__21501\,
            I => \N__21472\
        );

    \I__5074\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21472\
        );

    \I__5073\ : InMux
    port map (
            O => \N__21499\,
            I => \N__21467\
        );

    \I__5072\ : InMux
    port map (
            O => \N__21498\,
            I => \N__21467\
        );

    \I__5071\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21464\
        );

    \I__5070\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21459\
        );

    \I__5069\ : InMux
    port map (
            O => \N__21495\,
            I => \N__21459\
        );

    \I__5068\ : Span4Mux_h
    port map (
            O => \N__21492\,
            I => \N__21456\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__21489\,
            I => \N__21453\
        );

    \I__5066\ : Span4Mux_v
    port map (
            O => \N__21484\,
            I => \N__21448\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__21481\,
            I => \N__21448\
        );

    \I__5064\ : InMux
    port map (
            O => \N__21480\,
            I => \N__21445\
        );

    \I__5063\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21442\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__21472\,
            I => \N__21437\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__21467\,
            I => \N__21437\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__21464\,
            I => \N__21432\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__21459\,
            I => \N__21432\
        );

    \I__5058\ : Odrv4
    port map (
            O => \N__21456\,
            I => \Lab_UT.scctrl.N_223\
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__21453\,
            I => \Lab_UT.scctrl.N_223\
        );

    \I__5056\ : Odrv4
    port map (
            O => \N__21448\,
            I => \Lab_UT.scctrl.N_223\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__21445\,
            I => \Lab_UT.scctrl.N_223\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__21442\,
            I => \Lab_UT.scctrl.N_223\
        );

    \I__5053\ : Odrv4
    port map (
            O => \N__21437\,
            I => \Lab_UT.scctrl.N_223\
        );

    \I__5052\ : Odrv12
    port map (
            O => \N__21432\,
            I => \Lab_UT.scctrl.N_223\
        );

    \I__5051\ : CascadeMux
    port map (
            O => \N__21417\,
            I => \N__21405\
        );

    \I__5050\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21399\
        );

    \I__5049\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21392\
        );

    \I__5048\ : InMux
    port map (
            O => \N__21414\,
            I => \N__21392\
        );

    \I__5047\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21392\
        );

    \I__5046\ : InMux
    port map (
            O => \N__21412\,
            I => \N__21381\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21381\
        );

    \I__5044\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21381\
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__21409\,
            I => \N__21378\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21374\
        );

    \I__5041\ : InMux
    port map (
            O => \N__21405\,
            I => \N__21371\
        );

    \I__5040\ : InMux
    port map (
            O => \N__21404\,
            I => \N__21366\
        );

    \I__5039\ : InMux
    port map (
            O => \N__21403\,
            I => \N__21359\
        );

    \I__5038\ : InMux
    port map (
            O => \N__21402\,
            I => \N__21359\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__21399\,
            I => \N__21356\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21353\
        );

    \I__5035\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21350\
        );

    \I__5034\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21347\
        );

    \I__5033\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21342\
        );

    \I__5032\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21342\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__21381\,
            I => \N__21339\
        );

    \I__5030\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21334\
        );

    \I__5029\ : InMux
    port map (
            O => \N__21377\,
            I => \N__21334\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__21374\,
            I => \N__21329\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__21371\,
            I => \N__21326\
        );

    \I__5026\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21321\
        );

    \I__5025\ : InMux
    port map (
            O => \N__21369\,
            I => \N__21321\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__21366\,
            I => \N__21318\
        );

    \I__5023\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21309\
        );

    \I__5022\ : InMux
    port map (
            O => \N__21364\,
            I => \N__21309\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__21359\,
            I => \N__21306\
        );

    \I__5020\ : Span4Mux_v
    port map (
            O => \N__21356\,
            I => \N__21300\
        );

    \I__5019\ : Span4Mux_v
    port map (
            O => \N__21353\,
            I => \N__21300\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__21350\,
            I => \N__21297\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__21347\,
            I => \N__21288\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__21342\,
            I => \N__21288\
        );

    \I__5015\ : Span4Mux_v
    port map (
            O => \N__21339\,
            I => \N__21288\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__21334\,
            I => \N__21288\
        );

    \I__5013\ : InMux
    port map (
            O => \N__21333\,
            I => \N__21283\
        );

    \I__5012\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21283\
        );

    \I__5011\ : Span4Mux_v
    port map (
            O => \N__21329\,
            I => \N__21280\
        );

    \I__5010\ : Span4Mux_v
    port map (
            O => \N__21326\,
            I => \N__21275\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__21321\,
            I => \N__21275\
        );

    \I__5008\ : Span4Mux_s2_h
    port map (
            O => \N__21318\,
            I => \N__21272\
        );

    \I__5007\ : InMux
    port map (
            O => \N__21317\,
            I => \N__21267\
        );

    \I__5006\ : InMux
    port map (
            O => \N__21316\,
            I => \N__21267\
        );

    \I__5005\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21264\
        );

    \I__5004\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21261\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__21309\,
            I => \N__21258\
        );

    \I__5002\ : Span4Mux_s3_h
    port map (
            O => \N__21306\,
            I => \N__21255\
        );

    \I__5001\ : InMux
    port map (
            O => \N__21305\,
            I => \N__21252\
        );

    \I__5000\ : Span4Mux_h
    port map (
            O => \N__21300\,
            I => \N__21243\
        );

    \I__4999\ : Span4Mux_h
    port map (
            O => \N__21297\,
            I => \N__21243\
        );

    \I__4998\ : Span4Mux_v
    port map (
            O => \N__21288\,
            I => \N__21243\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__21283\,
            I => \N__21243\
        );

    \I__4996\ : Span4Mux_v
    port map (
            O => \N__21280\,
            I => \N__21236\
        );

    \I__4995\ : Span4Mux_v
    port map (
            O => \N__21275\,
            I => \N__21236\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__21272\,
            I => \N__21236\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__21267\,
            I => \Lab_UT.scctrl.stateZ0Z_0\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__21264\,
            I => \Lab_UT.scctrl.stateZ0Z_0\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__21261\,
            I => \Lab_UT.scctrl.stateZ0Z_0\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__21258\,
            I => \Lab_UT.scctrl.stateZ0Z_0\
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__21255\,
            I => \Lab_UT.scctrl.stateZ0Z_0\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__21252\,
            I => \Lab_UT.scctrl.stateZ0Z_0\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__21243\,
            I => \Lab_UT.scctrl.stateZ0Z_0\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__21236\,
            I => \Lab_UT.scctrl.stateZ0Z_0\
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__21219\,
            I => \N__21216\
        );

    \I__4984\ : InMux
    port map (
            O => \N__21216\,
            I => \N__21213\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__21213\,
            I => \N__21210\
        );

    \I__4982\ : Span4Mux_v
    port map (
            O => \N__21210\,
            I => \N__21207\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__21207\,
            I => \Lab_UT.scctrl.N_5_0\
        );

    \I__4980\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21201\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__21201\,
            I => \N__21198\
        );

    \I__4978\ : Span4Mux_v
    port map (
            O => \N__21198\,
            I => \N__21195\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__21195\,
            I => \Lab_UT.scctrl.G_10_i_a7_0_2\
        );

    \I__4976\ : IoInMux
    port map (
            O => \N__21192\,
            I => \N__21189\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__21189\,
            I => \N__21184\
        );

    \I__4974\ : InMux
    port map (
            O => \N__21188\,
            I => \N__21181\
        );

    \I__4973\ : InMux
    port map (
            O => \N__21187\,
            I => \N__21178\
        );

    \I__4972\ : Span4Mux_s1_v
    port map (
            O => \N__21184\,
            I => \N__21175\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__21181\,
            I => \N__21172\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__21178\,
            I => \N__21169\
        );

    \I__4969\ : Span4Mux_v
    port map (
            O => \N__21175\,
            I => \N__21166\
        );

    \I__4968\ : Span4Mux_v
    port map (
            O => \N__21172\,
            I => \N__21161\
        );

    \I__4967\ : Span4Mux_s1_h
    port map (
            O => \N__21169\,
            I => \N__21161\
        );

    \I__4966\ : Span4Mux_h
    port map (
            O => \N__21166\,
            I => \N__21158\
        );

    \I__4965\ : Span4Mux_h
    port map (
            O => \N__21161\,
            I => \N__21155\
        );

    \I__4964\ : Odrv4
    port map (
            O => \N__21158\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__21155\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4962\ : ClkMux
    port map (
            O => \N__21150\,
            I => \N__20907\
        );

    \I__4961\ : ClkMux
    port map (
            O => \N__21149\,
            I => \N__20907\
        );

    \I__4960\ : ClkMux
    port map (
            O => \N__21148\,
            I => \N__20907\
        );

    \I__4959\ : ClkMux
    port map (
            O => \N__21147\,
            I => \N__20907\
        );

    \I__4958\ : ClkMux
    port map (
            O => \N__21146\,
            I => \N__20907\
        );

    \I__4957\ : ClkMux
    port map (
            O => \N__21145\,
            I => \N__20907\
        );

    \I__4956\ : ClkMux
    port map (
            O => \N__21144\,
            I => \N__20907\
        );

    \I__4955\ : ClkMux
    port map (
            O => \N__21143\,
            I => \N__20907\
        );

    \I__4954\ : ClkMux
    port map (
            O => \N__21142\,
            I => \N__20907\
        );

    \I__4953\ : ClkMux
    port map (
            O => \N__21141\,
            I => \N__20907\
        );

    \I__4952\ : ClkMux
    port map (
            O => \N__21140\,
            I => \N__20907\
        );

    \I__4951\ : ClkMux
    port map (
            O => \N__21139\,
            I => \N__20907\
        );

    \I__4950\ : ClkMux
    port map (
            O => \N__21138\,
            I => \N__20907\
        );

    \I__4949\ : ClkMux
    port map (
            O => \N__21137\,
            I => \N__20907\
        );

    \I__4948\ : ClkMux
    port map (
            O => \N__21136\,
            I => \N__20907\
        );

    \I__4947\ : ClkMux
    port map (
            O => \N__21135\,
            I => \N__20907\
        );

    \I__4946\ : ClkMux
    port map (
            O => \N__21134\,
            I => \N__20907\
        );

    \I__4945\ : ClkMux
    port map (
            O => \N__21133\,
            I => \N__20907\
        );

    \I__4944\ : ClkMux
    port map (
            O => \N__21132\,
            I => \N__20907\
        );

    \I__4943\ : ClkMux
    port map (
            O => \N__21131\,
            I => \N__20907\
        );

    \I__4942\ : ClkMux
    port map (
            O => \N__21130\,
            I => \N__20907\
        );

    \I__4941\ : ClkMux
    port map (
            O => \N__21129\,
            I => \N__20907\
        );

    \I__4940\ : ClkMux
    port map (
            O => \N__21128\,
            I => \N__20907\
        );

    \I__4939\ : ClkMux
    port map (
            O => \N__21127\,
            I => \N__20907\
        );

    \I__4938\ : ClkMux
    port map (
            O => \N__21126\,
            I => \N__20907\
        );

    \I__4937\ : ClkMux
    port map (
            O => \N__21125\,
            I => \N__20907\
        );

    \I__4936\ : ClkMux
    port map (
            O => \N__21124\,
            I => \N__20907\
        );

    \I__4935\ : ClkMux
    port map (
            O => \N__21123\,
            I => \N__20907\
        );

    \I__4934\ : ClkMux
    port map (
            O => \N__21122\,
            I => \N__20907\
        );

    \I__4933\ : ClkMux
    port map (
            O => \N__21121\,
            I => \N__20907\
        );

    \I__4932\ : ClkMux
    port map (
            O => \N__21120\,
            I => \N__20907\
        );

    \I__4931\ : ClkMux
    port map (
            O => \N__21119\,
            I => \N__20907\
        );

    \I__4930\ : ClkMux
    port map (
            O => \N__21118\,
            I => \N__20907\
        );

    \I__4929\ : ClkMux
    port map (
            O => \N__21117\,
            I => \N__20907\
        );

    \I__4928\ : ClkMux
    port map (
            O => \N__21116\,
            I => \N__20907\
        );

    \I__4927\ : ClkMux
    port map (
            O => \N__21115\,
            I => \N__20907\
        );

    \I__4926\ : ClkMux
    port map (
            O => \N__21114\,
            I => \N__20907\
        );

    \I__4925\ : ClkMux
    port map (
            O => \N__21113\,
            I => \N__20907\
        );

    \I__4924\ : ClkMux
    port map (
            O => \N__21112\,
            I => \N__20907\
        );

    \I__4923\ : ClkMux
    port map (
            O => \N__21111\,
            I => \N__20907\
        );

    \I__4922\ : ClkMux
    port map (
            O => \N__21110\,
            I => \N__20907\
        );

    \I__4921\ : ClkMux
    port map (
            O => \N__21109\,
            I => \N__20907\
        );

    \I__4920\ : ClkMux
    port map (
            O => \N__21108\,
            I => \N__20907\
        );

    \I__4919\ : ClkMux
    port map (
            O => \N__21107\,
            I => \N__20907\
        );

    \I__4918\ : ClkMux
    port map (
            O => \N__21106\,
            I => \N__20907\
        );

    \I__4917\ : ClkMux
    port map (
            O => \N__21105\,
            I => \N__20907\
        );

    \I__4916\ : ClkMux
    port map (
            O => \N__21104\,
            I => \N__20907\
        );

    \I__4915\ : ClkMux
    port map (
            O => \N__21103\,
            I => \N__20907\
        );

    \I__4914\ : ClkMux
    port map (
            O => \N__21102\,
            I => \N__20907\
        );

    \I__4913\ : ClkMux
    port map (
            O => \N__21101\,
            I => \N__20907\
        );

    \I__4912\ : ClkMux
    port map (
            O => \N__21100\,
            I => \N__20907\
        );

    \I__4911\ : ClkMux
    port map (
            O => \N__21099\,
            I => \N__20907\
        );

    \I__4910\ : ClkMux
    port map (
            O => \N__21098\,
            I => \N__20907\
        );

    \I__4909\ : ClkMux
    port map (
            O => \N__21097\,
            I => \N__20907\
        );

    \I__4908\ : ClkMux
    port map (
            O => \N__21096\,
            I => \N__20907\
        );

    \I__4907\ : ClkMux
    port map (
            O => \N__21095\,
            I => \N__20907\
        );

    \I__4906\ : ClkMux
    port map (
            O => \N__21094\,
            I => \N__20907\
        );

    \I__4905\ : ClkMux
    port map (
            O => \N__21093\,
            I => \N__20907\
        );

    \I__4904\ : ClkMux
    port map (
            O => \N__21092\,
            I => \N__20907\
        );

    \I__4903\ : ClkMux
    port map (
            O => \N__21091\,
            I => \N__20907\
        );

    \I__4902\ : ClkMux
    port map (
            O => \N__21090\,
            I => \N__20907\
        );

    \I__4901\ : ClkMux
    port map (
            O => \N__21089\,
            I => \N__20907\
        );

    \I__4900\ : ClkMux
    port map (
            O => \N__21088\,
            I => \N__20907\
        );

    \I__4899\ : ClkMux
    port map (
            O => \N__21087\,
            I => \N__20907\
        );

    \I__4898\ : ClkMux
    port map (
            O => \N__21086\,
            I => \N__20907\
        );

    \I__4897\ : ClkMux
    port map (
            O => \N__21085\,
            I => \N__20907\
        );

    \I__4896\ : ClkMux
    port map (
            O => \N__21084\,
            I => \N__20907\
        );

    \I__4895\ : ClkMux
    port map (
            O => \N__21083\,
            I => \N__20907\
        );

    \I__4894\ : ClkMux
    port map (
            O => \N__21082\,
            I => \N__20907\
        );

    \I__4893\ : ClkMux
    port map (
            O => \N__21081\,
            I => \N__20907\
        );

    \I__4892\ : ClkMux
    port map (
            O => \N__21080\,
            I => \N__20907\
        );

    \I__4891\ : ClkMux
    port map (
            O => \N__21079\,
            I => \N__20907\
        );

    \I__4890\ : ClkMux
    port map (
            O => \N__21078\,
            I => \N__20907\
        );

    \I__4889\ : ClkMux
    port map (
            O => \N__21077\,
            I => \N__20907\
        );

    \I__4888\ : ClkMux
    port map (
            O => \N__21076\,
            I => \N__20907\
        );

    \I__4887\ : ClkMux
    port map (
            O => \N__21075\,
            I => \N__20907\
        );

    \I__4886\ : ClkMux
    port map (
            O => \N__21074\,
            I => \N__20907\
        );

    \I__4885\ : ClkMux
    port map (
            O => \N__21073\,
            I => \N__20907\
        );

    \I__4884\ : ClkMux
    port map (
            O => \N__21072\,
            I => \N__20907\
        );

    \I__4883\ : ClkMux
    port map (
            O => \N__21071\,
            I => \N__20907\
        );

    \I__4882\ : ClkMux
    port map (
            O => \N__21070\,
            I => \N__20907\
        );

    \I__4881\ : GlobalMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__4880\ : gio2CtrlBuf
    port map (
            O => \N__20904\,
            I => clk_g
        );

    \I__4879\ : CEMux
    port map (
            O => \N__20901\,
            I => \N__20896\
        );

    \I__4878\ : CEMux
    port map (
            O => \N__20900\,
            I => \N__20893\
        );

    \I__4877\ : CEMux
    port map (
            O => \N__20899\,
            I => \N__20889\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__20896\,
            I => \N__20886\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__20893\,
            I => \N__20883\
        );

    \I__4874\ : CEMux
    port map (
            O => \N__20892\,
            I => \N__20880\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__20889\,
            I => \N__20877\
        );

    \I__4872\ : Span4Mux_h
    port map (
            O => \N__20886\,
            I => \N__20874\
        );

    \I__4871\ : Span4Mux_h
    port map (
            O => \N__20883\,
            I => \N__20869\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__20880\,
            I => \N__20869\
        );

    \I__4869\ : Odrv4
    port map (
            O => \N__20877\,
            I => \Lab_UT.scctrl.next_state_RNIN96CP1Z0Z_3\
        );

    \I__4868\ : Odrv4
    port map (
            O => \N__20874\,
            I => \Lab_UT.scctrl.next_state_RNIN96CP1Z0Z_3\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__20869\,
            I => \Lab_UT.scctrl.next_state_RNIN96CP1Z0Z_3\
        );

    \I__4866\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20859\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__20859\,
            I => \N__20804\
        );

    \I__4864\ : SRMux
    port map (
            O => \N__20858\,
            I => \N__20697\
        );

    \I__4863\ : SRMux
    port map (
            O => \N__20857\,
            I => \N__20697\
        );

    \I__4862\ : SRMux
    port map (
            O => \N__20856\,
            I => \N__20697\
        );

    \I__4861\ : SRMux
    port map (
            O => \N__20855\,
            I => \N__20697\
        );

    \I__4860\ : SRMux
    port map (
            O => \N__20854\,
            I => \N__20697\
        );

    \I__4859\ : SRMux
    port map (
            O => \N__20853\,
            I => \N__20697\
        );

    \I__4858\ : SRMux
    port map (
            O => \N__20852\,
            I => \N__20697\
        );

    \I__4857\ : SRMux
    port map (
            O => \N__20851\,
            I => \N__20697\
        );

    \I__4856\ : SRMux
    port map (
            O => \N__20850\,
            I => \N__20697\
        );

    \I__4855\ : SRMux
    port map (
            O => \N__20849\,
            I => \N__20697\
        );

    \I__4854\ : SRMux
    port map (
            O => \N__20848\,
            I => \N__20697\
        );

    \I__4853\ : SRMux
    port map (
            O => \N__20847\,
            I => \N__20697\
        );

    \I__4852\ : SRMux
    port map (
            O => \N__20846\,
            I => \N__20697\
        );

    \I__4851\ : SRMux
    port map (
            O => \N__20845\,
            I => \N__20697\
        );

    \I__4850\ : SRMux
    port map (
            O => \N__20844\,
            I => \N__20697\
        );

    \I__4849\ : SRMux
    port map (
            O => \N__20843\,
            I => \N__20697\
        );

    \I__4848\ : SRMux
    port map (
            O => \N__20842\,
            I => \N__20697\
        );

    \I__4847\ : SRMux
    port map (
            O => \N__20841\,
            I => \N__20697\
        );

    \I__4846\ : SRMux
    port map (
            O => \N__20840\,
            I => \N__20697\
        );

    \I__4845\ : SRMux
    port map (
            O => \N__20839\,
            I => \N__20697\
        );

    \I__4844\ : SRMux
    port map (
            O => \N__20838\,
            I => \N__20697\
        );

    \I__4843\ : SRMux
    port map (
            O => \N__20837\,
            I => \N__20697\
        );

    \I__4842\ : SRMux
    port map (
            O => \N__20836\,
            I => \N__20697\
        );

    \I__4841\ : SRMux
    port map (
            O => \N__20835\,
            I => \N__20697\
        );

    \I__4840\ : SRMux
    port map (
            O => \N__20834\,
            I => \N__20697\
        );

    \I__4839\ : SRMux
    port map (
            O => \N__20833\,
            I => \N__20697\
        );

    \I__4838\ : SRMux
    port map (
            O => \N__20832\,
            I => \N__20697\
        );

    \I__4837\ : SRMux
    port map (
            O => \N__20831\,
            I => \N__20697\
        );

    \I__4836\ : SRMux
    port map (
            O => \N__20830\,
            I => \N__20697\
        );

    \I__4835\ : SRMux
    port map (
            O => \N__20829\,
            I => \N__20697\
        );

    \I__4834\ : SRMux
    port map (
            O => \N__20828\,
            I => \N__20697\
        );

    \I__4833\ : SRMux
    port map (
            O => \N__20827\,
            I => \N__20697\
        );

    \I__4832\ : SRMux
    port map (
            O => \N__20826\,
            I => \N__20697\
        );

    \I__4831\ : SRMux
    port map (
            O => \N__20825\,
            I => \N__20697\
        );

    \I__4830\ : SRMux
    port map (
            O => \N__20824\,
            I => \N__20697\
        );

    \I__4829\ : SRMux
    port map (
            O => \N__20823\,
            I => \N__20697\
        );

    \I__4828\ : SRMux
    port map (
            O => \N__20822\,
            I => \N__20697\
        );

    \I__4827\ : SRMux
    port map (
            O => \N__20821\,
            I => \N__20697\
        );

    \I__4826\ : SRMux
    port map (
            O => \N__20820\,
            I => \N__20697\
        );

    \I__4825\ : SRMux
    port map (
            O => \N__20819\,
            I => \N__20697\
        );

    \I__4824\ : SRMux
    port map (
            O => \N__20818\,
            I => \N__20697\
        );

    \I__4823\ : SRMux
    port map (
            O => \N__20817\,
            I => \N__20697\
        );

    \I__4822\ : SRMux
    port map (
            O => \N__20816\,
            I => \N__20697\
        );

    \I__4821\ : SRMux
    port map (
            O => \N__20815\,
            I => \N__20697\
        );

    \I__4820\ : SRMux
    port map (
            O => \N__20814\,
            I => \N__20697\
        );

    \I__4819\ : SRMux
    port map (
            O => \N__20813\,
            I => \N__20697\
        );

    \I__4818\ : SRMux
    port map (
            O => \N__20812\,
            I => \N__20697\
        );

    \I__4817\ : SRMux
    port map (
            O => \N__20811\,
            I => \N__20697\
        );

    \I__4816\ : SRMux
    port map (
            O => \N__20810\,
            I => \N__20697\
        );

    \I__4815\ : SRMux
    port map (
            O => \N__20809\,
            I => \N__20697\
        );

    \I__4814\ : SRMux
    port map (
            O => \N__20808\,
            I => \N__20697\
        );

    \I__4813\ : SRMux
    port map (
            O => \N__20807\,
            I => \N__20697\
        );

    \I__4812\ : Glb2LocalMux
    port map (
            O => \N__20804\,
            I => \N__20697\
        );

    \I__4811\ : GlobalMux
    port map (
            O => \N__20697\,
            I => \N__20694\
        );

    \I__4810\ : gio2CtrlBuf
    port map (
            O => \N__20694\,
            I => \resetGen_rst_1_iso_g\
        );

    \I__4809\ : CascadeMux
    port map (
            O => \N__20691\,
            I => \N__20687\
        );

    \I__4808\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20681\
        );

    \I__4807\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20681\
        );

    \I__4806\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20678\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__20681\,
            I => \N__20675\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__20678\,
            I => \N__20672\
        );

    \I__4803\ : Span4Mux_v
    port map (
            O => \N__20675\,
            I => \N__20669\
        );

    \I__4802\ : Odrv4
    port map (
            O => \N__20672\,
            I => \Lab_UT.scctrl.N_260\
        );

    \I__4801\ : Odrv4
    port map (
            O => \N__20669\,
            I => \Lab_UT.scctrl.N_260\
        );

    \I__4800\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20658\
        );

    \I__4799\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20652\
        );

    \I__4798\ : CascadeMux
    port map (
            O => \N__20662\,
            I => \N__20648\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__20661\,
            I => \N__20644\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__20658\,
            I => \N__20638\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20635\
        );

    \I__4794\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20632\
        );

    \I__4793\ : InMux
    port map (
            O => \N__20655\,
            I => \N__20629\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__20652\,
            I => \N__20626\
        );

    \I__4791\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20623\
        );

    \I__4790\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20620\
        );

    \I__4789\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20617\
        );

    \I__4788\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20614\
        );

    \I__4787\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20609\
        );

    \I__4786\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20609\
        );

    \I__4785\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20606\
        );

    \I__4784\ : Span4Mux_h
    port map (
            O => \N__20638\,
            I => \N__20596\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__20635\,
            I => \N__20596\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__20632\,
            I => \N__20596\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__20629\,
            I => \N__20596\
        );

    \I__4780\ : Span4Mux_h
    port map (
            O => \N__20626\,
            I => \N__20591\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__20623\,
            I => \N__20591\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__20620\,
            I => \N__20586\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__20617\,
            I => \N__20586\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__20614\,
            I => \N__20578\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20578\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__20606\,
            I => \N__20578\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__20605\,
            I => \N__20574\
        );

    \I__4772\ : Sp12to4
    port map (
            O => \N__20596\,
            I => \N__20571\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__20591\,
            I => \N__20566\
        );

    \I__4770\ : Span4Mux_v
    port map (
            O => \N__20586\,
            I => \N__20566\
        );

    \I__4769\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20563\
        );

    \I__4768\ : Span4Mux_h
    port map (
            O => \N__20578\,
            I => \N__20560\
        );

    \I__4767\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20557\
        );

    \I__4766\ : InMux
    port map (
            O => \N__20574\,
            I => \N__20554\
        );

    \I__4765\ : Odrv12
    port map (
            O => \N__20571\,
            I => \Lab_UT.scctrl.N_235\
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__20566\,
            I => \Lab_UT.scctrl.N_235\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__20563\,
            I => \Lab_UT.scctrl.N_235\
        );

    \I__4762\ : Odrv4
    port map (
            O => \N__20560\,
            I => \Lab_UT.scctrl.N_235\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__20557\,
            I => \Lab_UT.scctrl.N_235\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__20554\,
            I => \Lab_UT.scctrl.N_235\
        );

    \I__4759\ : IoInMux
    port map (
            O => \N__20541\,
            I => \N__20538\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__20538\,
            I => \N__20535\
        );

    \I__4757\ : IoSpan4Mux
    port map (
            O => \N__20535\,
            I => \N__20532\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__20532\,
            I => \N_55_i\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__20529\,
            I => \N__20525\
        );

    \I__4754\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20517\
        );

    \I__4753\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20514\
        );

    \I__4752\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20509\
        );

    \I__4751\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20505\
        );

    \I__4750\ : InMux
    port map (
            O => \N__20522\,
            I => \N__20502\
        );

    \I__4749\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20499\
        );

    \I__4748\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20496\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__20517\,
            I => \N__20491\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__20514\,
            I => \N__20491\
        );

    \I__4745\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20486\
        );

    \I__4744\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20486\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__20509\,
            I => \N__20483\
        );

    \I__4742\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20480\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20475\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__20502\,
            I => \N__20475\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__20499\,
            I => \N__20472\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__20496\,
            I => \Lab_UT.scctrl.state_i_1_0_rep1\
        );

    \I__4737\ : Odrv4
    port map (
            O => \N__20491\,
            I => \Lab_UT.scctrl.state_i_1_0_rep1\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__20486\,
            I => \Lab_UT.scctrl.state_i_1_0_rep1\
        );

    \I__4735\ : Odrv12
    port map (
            O => \N__20483\,
            I => \Lab_UT.scctrl.state_i_1_0_rep1\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__20480\,
            I => \Lab_UT.scctrl.state_i_1_0_rep1\
        );

    \I__4733\ : Odrv4
    port map (
            O => \N__20475\,
            I => \Lab_UT.scctrl.state_i_1_0_rep1\
        );

    \I__4732\ : Odrv4
    port map (
            O => \N__20472\,
            I => \Lab_UT.scctrl.state_i_1_0_rep1\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__20457\,
            I => \N__20453\
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__20456\,
            I => \N__20448\
        );

    \I__4729\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20444\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20452\,
            I => \N__20441\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20451\,
            I => \N__20438\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20448\,
            I => \N__20435\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__20447\,
            I => \N__20430\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__20444\,
            I => \N__20427\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__20441\,
            I => \N__20424\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__20438\,
            I => \N__20419\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__20435\,
            I => \N__20419\
        );

    \I__4720\ : InMux
    port map (
            O => \N__20434\,
            I => \N__20414\
        );

    \I__4719\ : InMux
    port map (
            O => \N__20433\,
            I => \N__20414\
        );

    \I__4718\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20411\
        );

    \I__4717\ : Span4Mux_h
    port map (
            O => \N__20427\,
            I => \N__20404\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__20424\,
            I => \N__20404\
        );

    \I__4715\ : Span4Mux_v
    port map (
            O => \N__20419\,
            I => \N__20404\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__20414\,
            I => \N__20399\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__20411\,
            I => \N__20399\
        );

    \I__4712\ : Span4Mux_v
    port map (
            O => \N__20404\,
            I => \N__20394\
        );

    \I__4711\ : Span4Mux_v
    port map (
            O => \N__20399\,
            I => \N__20394\
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__20394\,
            I => \Lab_UT.scctrl.state_2_rep1\
        );

    \I__4709\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20388\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__20388\,
            I => \Lab_UT.scctrl.N_13_1\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__20385\,
            I => \Lab_UT.scctrl.G_10_i_1_cascade_\
        );

    \I__4706\ : InMux
    port map (
            O => \N__20382\,
            I => \N__20379\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__20379\,
            I => \N__20376\
        );

    \I__4704\ : Span4Mux_s2_h
    port map (
            O => \N__20376\,
            I => \N__20372\
        );

    \I__4703\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20369\
        );

    \I__4702\ : Span4Mux_v
    port map (
            O => \N__20372\,
            I => \N__20366\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__20369\,
            I => \N__20363\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__20366\,
            I => \Lab_UT.scctrl.state_fast_2\
        );

    \I__4699\ : Odrv12
    port map (
            O => \N__20363\,
            I => \Lab_UT.scctrl.state_fast_2\
        );

    \I__4698\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20355\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__20355\,
            I => \N__20351\
        );

    \I__4696\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20347\
        );

    \I__4695\ : Span4Mux_s3_h
    port map (
            O => \N__20351\,
            I => \N__20344\
        );

    \I__4694\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20341\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__20347\,
            I => \N__20338\
        );

    \I__4692\ : Odrv4
    port map (
            O => \N__20344\,
            I => \Lab_UT.scctrl.state_i_1_fast_0\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__20341\,
            I => \Lab_UT.scctrl.state_i_1_fast_0\
        );

    \I__4690\ : Odrv12
    port map (
            O => \N__20338\,
            I => \Lab_UT.scctrl.state_i_1_fast_0\
        );

    \I__4689\ : CascadeMux
    port map (
            O => \N__20331\,
            I => \Lab_UT.scctrl.next_state_1_0_cascade_\
        );

    \I__4688\ : CascadeMux
    port map (
            O => \N__20328\,
            I => \N__20325\
        );

    \I__4687\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20322\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__20322\,
            I => \N__20319\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__20319\,
            I => \N__20316\
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__20316\,
            I => \Lab_UT.scctrl.N_356_1_0\
        );

    \I__4683\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20310\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__20310\,
            I => \N__20307\
        );

    \I__4681\ : Span4Mux_h
    port map (
            O => \N__20307\,
            I => \N__20304\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__20304\,
            I => \Lab_UT.scctrl.g0_9_a2_1\
        );

    \I__4679\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20298\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__20298\,
            I => \N__20295\
        );

    \I__4677\ : Span4Mux_s3_h
    port map (
            O => \N__20295\,
            I => \N__20292\
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__20292\,
            I => \Lab_UT.scctrl.g0_2_3_1\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__20289\,
            I => \N__20280\
        );

    \I__4674\ : CascadeMux
    port map (
            O => \N__20288\,
            I => \N__20277\
        );

    \I__4673\ : CascadeMux
    port map (
            O => \N__20287\,
            I => \N__20273\
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__20286\,
            I => \N__20270\
        );

    \I__4671\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20262\
        );

    \I__4670\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20262\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__20283\,
            I => \N__20259\
        );

    \I__4668\ : InMux
    port map (
            O => \N__20280\,
            I => \N__20253\
        );

    \I__4667\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20253\
        );

    \I__4666\ : InMux
    port map (
            O => \N__20276\,
            I => \N__20247\
        );

    \I__4665\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20236\
        );

    \I__4664\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20236\
        );

    \I__4663\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20236\
        );

    \I__4662\ : InMux
    port map (
            O => \N__20268\,
            I => \N__20236\
        );

    \I__4661\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20236\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20262\,
            I => \N__20233\
        );

    \I__4659\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20228\
        );

    \I__4658\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20228\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__20253\,
            I => \N__20225\
        );

    \I__4656\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20218\
        );

    \I__4655\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20218\
        );

    \I__4654\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20218\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__20247\,
            I => \N__20209\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__20236\,
            I => \N__20209\
        );

    \I__4651\ : Span4Mux_v
    port map (
            O => \N__20233\,
            I => \N__20209\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__20228\,
            I => \N__20209\
        );

    \I__4649\ : Span4Mux_v
    port map (
            O => \N__20225\,
            I => \N__20204\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__20218\,
            I => \N__20204\
        );

    \I__4647\ : Span4Mux_v
    port map (
            O => \N__20209\,
            I => \N__20199\
        );

    \I__4646\ : Span4Mux_h
    port map (
            O => \N__20204\,
            I => \N__20199\
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__20199\,
            I => \Lab_UT.scctrl.next_stateZ0Z_0\
        );

    \I__4644\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20193\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__4642\ : Span4Mux_h
    port map (
            O => \N__20190\,
            I => \N__20187\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__20187\,
            I => \Lab_UT.scctrl.g0_2_2_1\
        );

    \I__4640\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20172\
        );

    \I__4639\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20169\
        );

    \I__4638\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20166\
        );

    \I__4637\ : InMux
    port map (
            O => \N__20181\,
            I => \N__20161\
        );

    \I__4636\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20161\
        );

    \I__4635\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20158\
        );

    \I__4634\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20151\
        );

    \I__4633\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20151\
        );

    \I__4632\ : InMux
    port map (
            O => \N__20176\,
            I => \N__20151\
        );

    \I__4631\ : InMux
    port map (
            O => \N__20175\,
            I => \N__20148\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__20172\,
            I => \N__20145\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__20169\,
            I => \N__20142\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__20166\,
            I => \N__20136\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__20161\,
            I => \N__20131\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__20158\,
            I => \N__20131\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__20151\,
            I => \N__20128\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__20148\,
            I => \N__20125\
        );

    \I__4623\ : Span4Mux_v
    port map (
            O => \N__20145\,
            I => \N__20122\
        );

    \I__4622\ : Span4Mux_h
    port map (
            O => \N__20142\,
            I => \N__20119\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__20141\,
            I => \N__20115\
        );

    \I__4620\ : InMux
    port map (
            O => \N__20140\,
            I => \N__20111\
        );

    \I__4619\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20108\
        );

    \I__4618\ : Span4Mux_v
    port map (
            O => \N__20136\,
            I => \N__20103\
        );

    \I__4617\ : Span4Mux_v
    port map (
            O => \N__20131\,
            I => \N__20103\
        );

    \I__4616\ : Span4Mux_h
    port map (
            O => \N__20128\,
            I => \N__20100\
        );

    \I__4615\ : Span4Mux_v
    port map (
            O => \N__20125\,
            I => \N__20097\
        );

    \I__4614\ : Span4Mux_h
    port map (
            O => \N__20122\,
            I => \N__20092\
        );

    \I__4613\ : Span4Mux_v
    port map (
            O => \N__20119\,
            I => \N__20092\
        );

    \I__4612\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20089\
        );

    \I__4611\ : InMux
    port map (
            O => \N__20115\,
            I => \N__20084\
        );

    \I__4610\ : InMux
    port map (
            O => \N__20114\,
            I => \N__20084\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__20111\,
            I => \N__20079\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__20108\,
            I => \N__20079\
        );

    \I__4607\ : Span4Mux_h
    port map (
            O => \N__20103\,
            I => \N__20076\
        );

    \I__4606\ : Odrv4
    port map (
            O => \N__20100\,
            I => rst
        );

    \I__4605\ : Odrv4
    port map (
            O => \N__20097\,
            I => rst
        );

    \I__4604\ : Odrv4
    port map (
            O => \N__20092\,
            I => rst
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__20089\,
            I => rst
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__20084\,
            I => rst
        );

    \I__4601\ : Odrv12
    port map (
            O => \N__20079\,
            I => rst
        );

    \I__4600\ : Odrv4
    port map (
            O => \N__20076\,
            I => rst
        );

    \I__4599\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20058\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__20058\,
            I => \Lab_UT.scctrl.next_state_3_0\
        );

    \I__4597\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20049\
        );

    \I__4596\ : InMux
    port map (
            O => \N__20054\,
            I => \N__20046\
        );

    \I__4595\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20040\
        );

    \I__4594\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20040\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__20049\,
            I => \N__20034\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__20046\,
            I => \N__20031\
        );

    \I__4591\ : InMux
    port map (
            O => \N__20045\,
            I => \N__20028\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__20040\,
            I => \N__20025\
        );

    \I__4589\ : InMux
    port map (
            O => \N__20039\,
            I => \N__20018\
        );

    \I__4588\ : InMux
    port map (
            O => \N__20038\,
            I => \N__20018\
        );

    \I__4587\ : InMux
    port map (
            O => \N__20037\,
            I => \N__20018\
        );

    \I__4586\ : Span4Mux_s3_h
    port map (
            O => \N__20034\,
            I => \N__20011\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__20031\,
            I => \N__20006\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__20028\,
            I => \N__20006\
        );

    \I__4583\ : Span4Mux_h
    port map (
            O => \N__20025\,
            I => \N__20001\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__20018\,
            I => \N__20001\
        );

    \I__4581\ : InMux
    port map (
            O => \N__20017\,
            I => \N__19998\
        );

    \I__4580\ : InMux
    port map (
            O => \N__20016\,
            I => \N__19991\
        );

    \I__4579\ : InMux
    port map (
            O => \N__20015\,
            I => \N__19991\
        );

    \I__4578\ : InMux
    port map (
            O => \N__20014\,
            I => \N__19991\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__20011\,
            I => \Lab_UT.scctrl.next_stateZ0Z_1\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__20006\,
            I => \Lab_UT.scctrl.next_stateZ0Z_1\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__20001\,
            I => \Lab_UT.scctrl.next_stateZ0Z_1\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__19998\,
            I => \Lab_UT.scctrl.next_stateZ0Z_1\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__19991\,
            I => \Lab_UT.scctrl.next_stateZ0Z_1\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__19980\,
            I => \Lab_UT.scctrl.next_state_1_i_i_a2_1_0_1_cascade_\
        );

    \I__4571\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19973\
        );

    \I__4570\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19970\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__19973\,
            I => \N__19967\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__19970\,
            I => \N__19964\
        );

    \I__4567\ : Span4Mux_v
    port map (
            O => \N__19967\,
            I => \N__19959\
        );

    \I__4566\ : Span4Mux_v
    port map (
            O => \N__19964\,
            I => \N__19959\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__19959\,
            I => \Lab_UT.scctrl.next_state_rst_0_6\
        );

    \I__4564\ : InMux
    port map (
            O => \N__19956\,
            I => \N__19953\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__19953\,
            I => \N__19950\
        );

    \I__4562\ : Odrv12
    port map (
            O => \N__19950\,
            I => \Lab_UT.scctrl.N_398\
        );

    \I__4561\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19936\
        );

    \I__4560\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19936\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__19945\,
            I => \N__19931\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__19944\,
            I => \N__19927\
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__19943\,
            I => \N__19923\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__19942\,
            I => \N__19920\
        );

    \I__4555\ : CascadeMux
    port map (
            O => \N__19941\,
            I => \N__19917\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__19936\,
            I => \N__19914\
        );

    \I__4553\ : InMux
    port map (
            O => \N__19935\,
            I => \N__19911\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__19934\,
            I => \N__19908\
        );

    \I__4551\ : InMux
    port map (
            O => \N__19931\,
            I => \N__19903\
        );

    \I__4550\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19900\
        );

    \I__4549\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19891\
        );

    \I__4548\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19891\
        );

    \I__4547\ : InMux
    port map (
            O => \N__19923\,
            I => \N__19891\
        );

    \I__4546\ : InMux
    port map (
            O => \N__19920\,
            I => \N__19891\
        );

    \I__4545\ : InMux
    port map (
            O => \N__19917\,
            I => \N__19887\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__19914\,
            I => \N__19882\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__19911\,
            I => \N__19882\
        );

    \I__4542\ : InMux
    port map (
            O => \N__19908\,
            I => \N__19877\
        );

    \I__4541\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19877\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__19906\,
            I => \N__19874\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__19903\,
            I => \N__19870\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__19900\,
            I => \N__19865\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__19891\,
            I => \N__19865\
        );

    \I__4536\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19862\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__19887\,
            I => \N__19859\
        );

    \I__4534\ : Span4Mux_v
    port map (
            O => \N__19882\,
            I => \N__19854\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19854\
        );

    \I__4532\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19851\
        );

    \I__4531\ : CascadeMux
    port map (
            O => \N__19873\,
            I => \N__19848\
        );

    \I__4530\ : Span4Mux_v
    port map (
            O => \N__19870\,
            I => \N__19836\
        );

    \I__4529\ : Span4Mux_h
    port map (
            O => \N__19865\,
            I => \N__19836\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__19862\,
            I => \N__19836\
        );

    \I__4527\ : Span4Mux_v
    port map (
            O => \N__19859\,
            I => \N__19836\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__19854\,
            I => \N__19836\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__19851\,
            I => \N__19833\
        );

    \I__4524\ : InMux
    port map (
            O => \N__19848\,
            I => \N__19828\
        );

    \I__4523\ : InMux
    port map (
            O => \N__19847\,
            I => \N__19828\
        );

    \I__4522\ : Span4Mux_v
    port map (
            O => \N__19836\,
            I => \N__19825\
        );

    \I__4521\ : Span12Mux_s5_v
    port map (
            O => \N__19833\,
            I => \N__19822\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__19828\,
            I => \Lab_UT.scctrl.N_235_i_0\
        );

    \I__4519\ : Odrv4
    port map (
            O => \N__19825\,
            I => \Lab_UT.scctrl.N_235_i_0\
        );

    \I__4518\ : Odrv12
    port map (
            O => \N__19822\,
            I => \Lab_UT.scctrl.N_235_i_0\
        );

    \I__4517\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19810\
        );

    \I__4516\ : InMux
    port map (
            O => \N__19814\,
            I => \N__19807\
        );

    \I__4515\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19804\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__19810\,
            I => \N__19801\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__19807\,
            I => \N__19796\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__19804\,
            I => \N__19796\
        );

    \I__4511\ : Span4Mux_s3_h
    port map (
            O => \N__19801\,
            I => \N__19793\
        );

    \I__4510\ : Odrv12
    port map (
            O => \N__19796\,
            I => \Lab_UT.scctrl.N_240\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__19793\,
            I => \Lab_UT.scctrl.N_240\
        );

    \I__4508\ : CascadeMux
    port map (
            O => \N__19788\,
            I => \N__19785\
        );

    \I__4507\ : InMux
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__19782\,
            I => \N__19779\
        );

    \I__4505\ : Span4Mux_s2_h
    port map (
            O => \N__19779\,
            I => \N__19776\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__19776\,
            I => \N__19773\
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__19773\,
            I => \Lab_UT.scctrl.N_296\
        );

    \I__4502\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19767\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19767\,
            I => \N__19764\
        );

    \I__4500\ : Odrv12
    port map (
            O => \N__19764\,
            I => \Lab_UT.scctrl.state_1_ret_1_RNICEVZ0Z81\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__19761\,
            I => \Lab_UT.scctrl.G_24_i_1_cascade_\
        );

    \I__4498\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__19755\,
            I => \N__19752\
        );

    \I__4496\ : Odrv12
    port map (
            O => \N__19752\,
            I => \Lab_UT.scctrl.N_13_2\
        );

    \I__4495\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19745\
        );

    \I__4494\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19742\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__19745\,
            I => \N__19737\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__19742\,
            I => \N__19737\
        );

    \I__4491\ : Span4Mux_h
    port map (
            O => \N__19737\,
            I => \N__19734\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__19734\,
            I => \Lab_UT.scctrl.rst_retZ0\
        );

    \I__4489\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19722\
        );

    \I__4488\ : CascadeMux
    port map (
            O => \N__19730\,
            I => \N__19719\
        );

    \I__4487\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19716\
        );

    \I__4486\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19713\
        );

    \I__4485\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19709\
        );

    \I__4484\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19706\
        );

    \I__4483\ : InMux
    port map (
            O => \N__19725\,
            I => \N__19703\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__19722\,
            I => \N__19700\
        );

    \I__4481\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19697\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__19716\,
            I => \N__19694\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__19713\,
            I => \N__19691\
        );

    \I__4478\ : InMux
    port map (
            O => \N__19712\,
            I => \N__19688\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__19709\,
            I => \N__19682\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__19706\,
            I => \N__19682\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__19703\,
            I => \N__19676\
        );

    \I__4474\ : Span4Mux_v
    port map (
            O => \N__19700\,
            I => \N__19676\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__19697\,
            I => \N__19671\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__19694\,
            I => \N__19671\
        );

    \I__4471\ : Span4Mux_h
    port map (
            O => \N__19691\,
            I => \N__19664\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__19688\,
            I => \N__19664\
        );

    \I__4469\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19661\
        );

    \I__4468\ : Span4Mux_s2_h
    port map (
            O => \N__19682\,
            I => \N__19658\
        );

    \I__4467\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19655\
        );

    \I__4466\ : Span4Mux_h
    port map (
            O => \N__19676\,
            I => \N__19650\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__19671\,
            I => \N__19650\
        );

    \I__4464\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19645\
        );

    \I__4463\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19645\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__19664\,
            I => \Lab_UT.scctrl.state_i_2_2\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__19661\,
            I => \Lab_UT.scctrl.state_i_2_2\
        );

    \I__4460\ : Odrv4
    port map (
            O => \N__19658\,
            I => \Lab_UT.scctrl.state_i_2_2\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__19655\,
            I => \Lab_UT.scctrl.state_i_2_2\
        );

    \I__4458\ : Odrv4
    port map (
            O => \N__19650\,
            I => \Lab_UT.scctrl.state_i_2_2\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__19645\,
            I => \Lab_UT.scctrl.state_i_2_2\
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__19632\,
            I => \Lab_UT.scctrl.N_12_cascade_\
        );

    \I__4455\ : InMux
    port map (
            O => \N__19629\,
            I => \N__19626\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__19626\,
            I => \N__19623\
        );

    \I__4453\ : Odrv12
    port map (
            O => \N__19623\,
            I => \Lab_UT.scctrl.N_8_0\
        );

    \I__4452\ : InMux
    port map (
            O => \N__19620\,
            I => \N__19617\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__19617\,
            I => \N__19614\
        );

    \I__4450\ : Span4Mux_h
    port map (
            O => \N__19614\,
            I => \N__19611\
        );

    \I__4449\ : Odrv4
    port map (
            O => \N__19611\,
            I => \Lab_UT.scctrl.g0_9_a2_4\
        );

    \I__4448\ : CascadeMux
    port map (
            O => \N__19608\,
            I => \N__19604\
        );

    \I__4447\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19600\
        );

    \I__4446\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19591\
        );

    \I__4445\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19591\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__19600\,
            I => \N__19588\
        );

    \I__4443\ : InMux
    port map (
            O => \N__19599\,
            I => \N__19581\
        );

    \I__4442\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19581\
        );

    \I__4441\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19581\
        );

    \I__4440\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19578\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__19591\,
            I => \N__19574\
        );

    \I__4438\ : Span4Mux_v
    port map (
            O => \N__19588\,
            I => \N__19567\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__19581\,
            I => \N__19567\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__19578\,
            I => \N__19564\
        );

    \I__4435\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19561\
        );

    \I__4434\ : Span4Mux_h
    port map (
            O => \N__19574\,
            I => \N__19558\
        );

    \I__4433\ : InMux
    port map (
            O => \N__19573\,
            I => \N__19553\
        );

    \I__4432\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19553\
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__19567\,
            I => \Lab_UT.scctrl.state_3_rep1\
        );

    \I__4430\ : Odrv4
    port map (
            O => \N__19564\,
            I => \Lab_UT.scctrl.state_3_rep1\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__19561\,
            I => \Lab_UT.scctrl.state_3_rep1\
        );

    \I__4428\ : Odrv4
    port map (
            O => \N__19558\,
            I => \Lab_UT.scctrl.state_3_rep1\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__19553\,
            I => \Lab_UT.scctrl.state_3_rep1\
        );

    \I__4426\ : InMux
    port map (
            O => \N__19542\,
            I => \N__19539\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__19539\,
            I => \Lab_UT.scctrl.g0_9_a3_0_0\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__19536\,
            I => \N__19531\
        );

    \I__4423\ : CascadeMux
    port map (
            O => \N__19535\,
            I => \N__19526\
        );

    \I__4422\ : CascadeMux
    port map (
            O => \N__19534\,
            I => \N__19522\
        );

    \I__4421\ : InMux
    port map (
            O => \N__19531\,
            I => \N__19513\
        );

    \I__4420\ : InMux
    port map (
            O => \N__19530\,
            I => \N__19513\
        );

    \I__4419\ : InMux
    port map (
            O => \N__19529\,
            I => \N__19500\
        );

    \I__4418\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19500\
        );

    \I__4417\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19500\
        );

    \I__4416\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19500\
        );

    \I__4415\ : InMux
    port map (
            O => \N__19521\,
            I => \N__19500\
        );

    \I__4414\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19500\
        );

    \I__4413\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19497\
        );

    \I__4412\ : InMux
    port map (
            O => \N__19518\,
            I => \N__19489\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__19513\,
            I => \N__19484\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__19500\,
            I => \N__19484\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__19497\,
            I => \N__19481\
        );

    \I__4408\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19476\
        );

    \I__4407\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19476\
        );

    \I__4406\ : InMux
    port map (
            O => \N__19494\,
            I => \N__19473\
        );

    \I__4405\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19470\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19492\,
            I => \N__19467\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19489\,
            I => \N__19464\
        );

    \I__4402\ : Span4Mux_v
    port map (
            O => \N__19484\,
            I => \N__19457\
        );

    \I__4401\ : Span4Mux_s3_h
    port map (
            O => \N__19481\,
            I => \N__19457\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__19476\,
            I => \N__19457\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__19473\,
            I => \N__19454\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__19470\,
            I => \N__19451\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__19467\,
            I => \N__19444\
        );

    \I__4396\ : Span4Mux_s3_h
    port map (
            O => \N__19464\,
            I => \N__19444\
        );

    \I__4395\ : Span4Mux_v
    port map (
            O => \N__19457\,
            I => \N__19444\
        );

    \I__4394\ : Span12Mux_s10_v
    port map (
            O => \N__19454\,
            I => \N__19441\
        );

    \I__4393\ : Odrv12
    port map (
            O => \N__19451\,
            I => \Lab_UT.scctrl.next_stateZ0Z_3\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__19444\,
            I => \Lab_UT.scctrl.next_stateZ0Z_3\
        );

    \I__4391\ : Odrv12
    port map (
            O => \N__19441\,
            I => \Lab_UT.scctrl.next_stateZ0Z_3\
        );

    \I__4390\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19430\
        );

    \I__4389\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19427\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__19430\,
            I => \N__19424\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__19427\,
            I => \N__19421\
        );

    \I__4386\ : Span4Mux_h
    port map (
            O => \N__19424\,
            I => \N__19418\
        );

    \I__4385\ : Span4Mux_s2_h
    port map (
            O => \N__19421\,
            I => \N__19415\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__19418\,
            I => \Lab_UT.scctrl.next_state_0_1\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__19415\,
            I => \Lab_UT.scctrl.next_state_0_1\
        );

    \I__4382\ : CascadeMux
    port map (
            O => \N__19410\,
            I => \Lab_UT.scctrl.m90_i_o6_0_0_cascade_\
        );

    \I__4381\ : InMux
    port map (
            O => \N__19407\,
            I => \N__19404\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__19404\,
            I => \N__19401\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__19401\,
            I => \N__19398\
        );

    \I__4378\ : Span4Mux_s1_h
    port map (
            O => \N__19398\,
            I => \N__19395\
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__19395\,
            I => \Lab_UT.scctrl.N_404_1\
        );

    \I__4376\ : InMux
    port map (
            O => \N__19392\,
            I => \N__19386\
        );

    \I__4375\ : InMux
    port map (
            O => \N__19391\,
            I => \N__19383\
        );

    \I__4374\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19380\
        );

    \I__4373\ : InMux
    port map (
            O => \N__19389\,
            I => \N__19377\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__19386\,
            I => \N__19373\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__19383\,
            I => \N__19370\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__19380\,
            I => \N__19366\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__19377\,
            I => \N__19363\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19360\
        );

    \I__4367\ : Span4Mux_v
    port map (
            O => \N__19373\,
            I => \N__19355\
        );

    \I__4366\ : Span4Mux_h
    port map (
            O => \N__19370\,
            I => \N__19355\
        );

    \I__4365\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19352\
        );

    \I__4364\ : Odrv12
    port map (
            O => \N__19366\,
            I => \Lab_UT.scctrl.N_401\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__19363\,
            I => \Lab_UT.scctrl.N_401\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__19360\,
            I => \Lab_UT.scctrl.N_401\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__19355\,
            I => \Lab_UT.scctrl.N_401\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__19352\,
            I => \Lab_UT.scctrl.N_401\
        );

    \I__4359\ : InMux
    port map (
            O => \N__19341\,
            I => \N__19337\
        );

    \I__4358\ : InMux
    port map (
            O => \N__19340\,
            I => \N__19334\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__19337\,
            I => \N__19328\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__19334\,
            I => \N__19325\
        );

    \I__4355\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19322\
        );

    \I__4354\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19317\
        );

    \I__4353\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19317\
        );

    \I__4352\ : Span4Mux_h
    port map (
            O => \N__19328\,
            I => \N__19312\
        );

    \I__4351\ : Span4Mux_h
    port map (
            O => \N__19325\,
            I => \N__19309\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__19322\,
            I => \N__19304\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__19317\,
            I => \N__19304\
        );

    \I__4348\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19301\
        );

    \I__4347\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19298\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__19312\,
            I => \Lab_UT.scctrl.N_399\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__19309\,
            I => \Lab_UT.scctrl.N_399\
        );

    \I__4344\ : Odrv12
    port map (
            O => \N__19304\,
            I => \Lab_UT.scctrl.N_399\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__19301\,
            I => \Lab_UT.scctrl.N_399\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__19298\,
            I => \Lab_UT.scctrl.N_399\
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__19287\,
            I => \Lab_UT.scctrl.g0_2_2_cascade_\
        );

    \I__4340\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19281\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__19281\,
            I => \N__19278\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__19278\,
            I => \N__19275\
        );

    \I__4337\ : Odrv4
    port map (
            O => \N__19275\,
            I => \Lab_UT.scctrl.g0_2_3\
        );

    \I__4336\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19269\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__19269\,
            I => \N__19265\
        );

    \I__4334\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19262\
        );

    \I__4333\ : Span4Mux_s2_h
    port map (
            O => \N__19265\,
            I => \N__19259\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__19262\,
            I => \N__19256\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__19259\,
            I => \Lab_UT.scctrl.g0_1_3\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__19256\,
            I => \Lab_UT.scctrl.g0_1_3\
        );

    \I__4329\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19248\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__19248\,
            I => \N__19238\
        );

    \I__4327\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19235\
        );

    \I__4326\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19222\
        );

    \I__4325\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19222\
        );

    \I__4324\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19222\
        );

    \I__4323\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19222\
        );

    \I__4322\ : InMux
    port map (
            O => \N__19242\,
            I => \N__19222\
        );

    \I__4321\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19222\
        );

    \I__4320\ : Odrv4
    port map (
            O => \N__19238\,
            I => \Lab_UT.scctrl.next_state_rst_2_2\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19235\,
            I => \Lab_UT.scctrl.next_state_rst_2_2\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__19222\,
            I => \Lab_UT.scctrl.next_state_rst_2_2\
        );

    \I__4317\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19212\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__19212\,
            I => \Lab_UT.scctrl.N_13\
        );

    \I__4315\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19206\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__19206\,
            I => \N__19203\
        );

    \I__4313\ : Span4Mux_v
    port map (
            O => \N__19203\,
            I => \N__19200\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__19200\,
            I => \N__19197\
        );

    \I__4311\ : Span4Mux_h
    port map (
            O => \N__19197\,
            I => \N__19194\
        );

    \I__4310\ : Odrv4
    port map (
            O => \N__19194\,
            I => \Lab_UT.scctrl.N_404_0\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__19191\,
            I => \Lab_UT.scctrl.N_5_3_cascade_\
        );

    \I__4308\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19185\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__19185\,
            I => \N__19182\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__19182\,
            I => \Lab_UT.scctrl.N_12_0\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__19179\,
            I => \N__19176\
        );

    \I__4304\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19173\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__19173\,
            I => \N__19170\
        );

    \I__4302\ : Span4Mux_s2_h
    port map (
            O => \N__19170\,
            I => \N__19167\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__19167\,
            I => \Lab_UT.scctrl.G_18_i_a9_0\
        );

    \I__4300\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19161\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__19161\,
            I => \Lab_UT.scctrl.N_14_0\
        );

    \I__4298\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19148\
        );

    \I__4297\ : CascadeMux
    port map (
            O => \N__19157\,
            I => \N__19145\
        );

    \I__4296\ : CascadeMux
    port map (
            O => \N__19156\,
            I => \N__19141\
        );

    \I__4295\ : InMux
    port map (
            O => \N__19155\,
            I => \N__19134\
        );

    \I__4294\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19134\
        );

    \I__4293\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19134\
        );

    \I__4292\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19126\
        );

    \I__4291\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19126\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__19148\,
            I => \N__19122\
        );

    \I__4289\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19117\
        );

    \I__4288\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19117\
        );

    \I__4287\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19114\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__19134\,
            I => \N__19111\
        );

    \I__4285\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19108\
        );

    \I__4284\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19105\
        );

    \I__4283\ : InMux
    port map (
            O => \N__19131\,
            I => \N__19100\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__19126\,
            I => \N__19097\
        );

    \I__4281\ : InMux
    port map (
            O => \N__19125\,
            I => \N__19094\
        );

    \I__4280\ : Span4Mux_v
    port map (
            O => \N__19122\,
            I => \N__19085\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__19117\,
            I => \N__19085\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__19114\,
            I => \N__19085\
        );

    \I__4277\ : Span4Mux_v
    port map (
            O => \N__19111\,
            I => \N__19085\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__19108\,
            I => \N__19082\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__19105\,
            I => \N__19079\
        );

    \I__4274\ : InMux
    port map (
            O => \N__19104\,
            I => \N__19074\
        );

    \I__4273\ : InMux
    port map (
            O => \N__19103\,
            I => \N__19074\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__19100\,
            I => \N__19071\
        );

    \I__4271\ : Span4Mux_v
    port map (
            O => \N__19097\,
            I => \N__19068\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__19094\,
            I => \N__19065\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__19085\,
            I => \N__19062\
        );

    \I__4268\ : Span4Mux_v
    port map (
            O => \N__19082\,
            I => \N__19059\
        );

    \I__4267\ : Sp12to4
    port map (
            O => \N__19079\,
            I => \N__19054\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__19074\,
            I => \N__19054\
        );

    \I__4265\ : Span4Mux_s3_v
    port map (
            O => \N__19071\,
            I => \N__19049\
        );

    \I__4264\ : Span4Mux_v
    port map (
            O => \N__19068\,
            I => \N__19049\
        );

    \I__4263\ : Span4Mux_v
    port map (
            O => \N__19065\,
            I => \N__19042\
        );

    \I__4262\ : Span4Mux_v
    port map (
            O => \N__19062\,
            I => \N__19042\
        );

    \I__4261\ : Span4Mux_s0_h
    port map (
            O => \N__19059\,
            I => \N__19042\
        );

    \I__4260\ : Odrv12
    port map (
            O => \N__19054\,
            I => \Lab_UT.scctrl.stateZ0Z_2\
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__19049\,
            I => \Lab_UT.scctrl.stateZ0Z_2\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__19042\,
            I => \Lab_UT.scctrl.stateZ0Z_2\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__19035\,
            I => \N__19032\
        );

    \I__4256\ : InMux
    port map (
            O => \N__19032\,
            I => \N__19028\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__19031\,
            I => \N__19025\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__19028\,
            I => \N__19022\
        );

    \I__4253\ : InMux
    port map (
            O => \N__19025\,
            I => \N__19019\
        );

    \I__4252\ : Span4Mux_s2_h
    port map (
            O => \N__19022\,
            I => \N__19016\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__19019\,
            I => \N__19013\
        );

    \I__4250\ : Odrv4
    port map (
            O => \N__19016\,
            I => \Lab_UT.scctrl.N_5\
        );

    \I__4249\ : Odrv4
    port map (
            O => \N__19013\,
            I => \Lab_UT.scctrl.N_5\
        );

    \I__4248\ : CascadeMux
    port map (
            O => \N__19008\,
            I => \N__19005\
        );

    \I__4247\ : InMux
    port map (
            O => \N__19005\,
            I => \N__19002\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__19002\,
            I => \N__18999\
        );

    \I__4245\ : Span4Mux_h
    port map (
            O => \N__18999\,
            I => \N__18996\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__18996\,
            I => \Lab_UT.scctrl.N_21_0\
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__18993\,
            I => \Lab_UT.scctrl.G_10_i_o7_0_cascade_\
        );

    \I__4242\ : InMux
    port map (
            O => \N__18990\,
            I => \N__18987\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__18987\,
            I => \N__18984\
        );

    \I__4240\ : Span4Mux_s3_h
    port map (
            O => \N__18984\,
            I => \N__18981\
        );

    \I__4239\ : Odrv4
    port map (
            O => \N__18981\,
            I => \Lab_UT.scctrl.G_24_i_a7_4_2\
        );

    \I__4238\ : InMux
    port map (
            O => \N__18978\,
            I => \N__18975\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__18975\,
            I => \Lab_UT.scctrl.G_18_i_a9_0_2\
        );

    \I__4236\ : InMux
    port map (
            O => \N__18972\,
            I => \N__18969\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__18969\,
            I => \N__18966\
        );

    \I__4234\ : Span4Mux_v
    port map (
            O => \N__18966\,
            I => \N__18963\
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__18963\,
            I => \Lab_UT.scctrl.G_18_i_1\
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__18960\,
            I => \Lab_UT.scctrl.G_18_i_2_cascade_\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__18957\,
            I => \Lab_UT.scctrl.G_18_i_4_cascade_\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__18954\,
            I => \N__18951\
        );

    \I__4229\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18948\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__18948\,
            I => \N__18945\
        );

    \I__4227\ : Span4Mux_h
    port map (
            O => \N__18945\,
            I => \N__18942\
        );

    \I__4226\ : Span4Mux_v
    port map (
            O => \N__18942\,
            I => \N__18939\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__18939\,
            I => \Lab_UT.scctrl.N_8_0_0\
        );

    \I__4224\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18933\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__18933\,
            I => \N__18930\
        );

    \I__4222\ : Span4Mux_s3_h
    port map (
            O => \N__18930\,
            I => \N__18927\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__18927\,
            I => \Lab_UT.scctrl.g0_2_3_0\
        );

    \I__4220\ : InMux
    port map (
            O => \N__18924\,
            I => \N__18921\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__18921\,
            I => \N__18918\
        );

    \I__4218\ : Span4Mux_h
    port map (
            O => \N__18918\,
            I => \N__18915\
        );

    \I__4217\ : Span4Mux_v
    port map (
            O => \N__18915\,
            I => \N__18912\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__18912\,
            I => \Lab_UT.scctrl.g0_2_2_0\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__18909\,
            I => \Lab_UT.scctrl.next_state_2_0_cascade_\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18906\,
            I => \N__18900\
        );

    \I__4213\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18894\
        );

    \I__4212\ : InMux
    port map (
            O => \N__18904\,
            I => \N__18891\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__18903\,
            I => \N__18888\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__18900\,
            I => \N__18884\
        );

    \I__4209\ : InMux
    port map (
            O => \N__18899\,
            I => \N__18879\
        );

    \I__4208\ : InMux
    port map (
            O => \N__18898\,
            I => \N__18879\
        );

    \I__4207\ : InMux
    port map (
            O => \N__18897\,
            I => \N__18876\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__18894\,
            I => \N__18873\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__18891\,
            I => \N__18870\
        );

    \I__4204\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18865\
        );

    \I__4203\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18865\
        );

    \I__4202\ : Span4Mux_v
    port map (
            O => \N__18884\,
            I => \N__18862\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__18879\,
            I => \N__18858\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__18876\,
            I => \N__18849\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__18873\,
            I => \N__18849\
        );

    \I__4198\ : Span4Mux_v
    port map (
            O => \N__18870\,
            I => \N__18849\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__18865\,
            I => \N__18849\
        );

    \I__4196\ : Span4Mux_v
    port map (
            O => \N__18862\,
            I => \N__18846\
        );

    \I__4195\ : InMux
    port map (
            O => \N__18861\,
            I => \N__18843\
        );

    \I__4194\ : Span4Mux_h
    port map (
            O => \N__18858\,
            I => \N__18838\
        );

    \I__4193\ : Span4Mux_h
    port map (
            O => \N__18849\,
            I => \N__18838\
        );

    \I__4192\ : Odrv4
    port map (
            O => \N__18846\,
            I => \Lab_UT.scctrl.N_260_i_0\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__18843\,
            I => \Lab_UT.scctrl.N_260_i_0\
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__18838\,
            I => \Lab_UT.scctrl.N_260_i_0\
        );

    \I__4189\ : CascadeMux
    port map (
            O => \N__18831\,
            I => \N__18828\
        );

    \I__4188\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18825\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__18825\,
            I => \N__18822\
        );

    \I__4186\ : Span4Mux_v
    port map (
            O => \N__18822\,
            I => \N__18819\
        );

    \I__4185\ : Span4Mux_h
    port map (
            O => \N__18819\,
            I => \N__18816\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__18816\,
            I => \Lab_UT.scctrl.N_404_4\
        );

    \I__4183\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18809\
        );

    \I__4182\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18805\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__18809\,
            I => \N__18800\
        );

    \I__4180\ : InMux
    port map (
            O => \N__18808\,
            I => \N__18797\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__18805\,
            I => \N__18794\
        );

    \I__4178\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18789\
        );

    \I__4177\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18789\
        );

    \I__4176\ : Span4Mux_h
    port map (
            O => \N__18800\,
            I => \N__18776\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__18797\,
            I => \N__18773\
        );

    \I__4174\ : Span4Mux_s3_h
    port map (
            O => \N__18794\,
            I => \N__18770\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__18789\,
            I => \N__18767\
        );

    \I__4172\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18764\
        );

    \I__4171\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18757\
        );

    \I__4170\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18757\
        );

    \I__4169\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18757\
        );

    \I__4168\ : InMux
    port map (
            O => \N__18784\,
            I => \N__18748\
        );

    \I__4167\ : InMux
    port map (
            O => \N__18783\,
            I => \N__18748\
        );

    \I__4166\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18748\
        );

    \I__4165\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18743\
        );

    \I__4164\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18743\
        );

    \I__4163\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18740\
        );

    \I__4162\ : Span4Mux_v
    port map (
            O => \N__18776\,
            I => \N__18731\
        );

    \I__4161\ : Span4Mux_h
    port map (
            O => \N__18773\,
            I => \N__18731\
        );

    \I__4160\ : Span4Mux_h
    port map (
            O => \N__18770\,
            I => \N__18731\
        );

    \I__4159\ : Span4Mux_h
    port map (
            O => \N__18767\,
            I => \N__18731\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__18764\,
            I => \N__18728\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__18757\,
            I => \N__18725\
        );

    \I__4156\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18722\
        );

    \I__4155\ : InMux
    port map (
            O => \N__18755\,
            I => \N__18719\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__18748\,
            I => bu_rx_data_5
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__18743\,
            I => bu_rx_data_5
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__18740\,
            I => bu_rx_data_5
        );

    \I__4151\ : Odrv4
    port map (
            O => \N__18731\,
            I => bu_rx_data_5
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__18728\,
            I => bu_rx_data_5
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__18725\,
            I => bu_rx_data_5
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__18722\,
            I => bu_rx_data_5
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__18719\,
            I => bu_rx_data_5
        );

    \I__4146\ : InMux
    port map (
            O => \N__18702\,
            I => \N__18699\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__18699\,
            I => \N__18696\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__18696\,
            I => \N__18693\
        );

    \I__4143\ : Odrv4
    port map (
            O => \N__18693\,
            I => \Lab_UT.scctrl.g0_1_1_1\
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__18690\,
            I => \N__18671\
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__18689\,
            I => \N__18661\
        );

    \I__4140\ : InMux
    port map (
            O => \N__18688\,
            I => \N__18655\
        );

    \I__4139\ : InMux
    port map (
            O => \N__18687\,
            I => \N__18652\
        );

    \I__4138\ : InMux
    port map (
            O => \N__18686\,
            I => \N__18647\
        );

    \I__4137\ : InMux
    port map (
            O => \N__18685\,
            I => \N__18647\
        );

    \I__4136\ : InMux
    port map (
            O => \N__18684\,
            I => \N__18642\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18683\,
            I => \N__18642\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18633\
        );

    \I__4133\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18633\
        );

    \I__4132\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18633\
        );

    \I__4131\ : InMux
    port map (
            O => \N__18679\,
            I => \N__18633\
        );

    \I__4130\ : InMux
    port map (
            O => \N__18678\,
            I => \N__18624\
        );

    \I__4129\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18624\
        );

    \I__4128\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18624\
        );

    \I__4127\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18624\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18606\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18606\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18606\
        );

    \I__4123\ : InMux
    port map (
            O => \N__18669\,
            I => \N__18606\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18668\,
            I => \N__18606\
        );

    \I__4121\ : InMux
    port map (
            O => \N__18667\,
            I => \N__18606\
        );

    \I__4120\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18606\
        );

    \I__4119\ : InMux
    port map (
            O => \N__18665\,
            I => \N__18606\
        );

    \I__4118\ : InMux
    port map (
            O => \N__18664\,
            I => \N__18595\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18661\,
            I => \N__18595\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18660\,
            I => \N__18595\
        );

    \I__4115\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18595\
        );

    \I__4114\ : InMux
    port map (
            O => \N__18658\,
            I => \N__18595\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__18655\,
            I => \N__18590\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__18652\,
            I => \N__18590\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__18647\,
            I => \N__18587\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__18642\,
            I => \N__18580\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__18633\,
            I => \N__18580\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__18624\,
            I => \N__18580\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__18623\,
            I => \N__18577\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18571\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18595\,
            I => \N__18566\
        );

    \I__4104\ : Span4Mux_s2_v
    port map (
            O => \N__18590\,
            I => \N__18566\
        );

    \I__4103\ : Span4Mux_v
    port map (
            O => \N__18587\,
            I => \N__18561\
        );

    \I__4102\ : Span4Mux_v
    port map (
            O => \N__18580\,
            I => \N__18561\
        );

    \I__4101\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18558\
        );

    \I__4100\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18551\
        );

    \I__4099\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18551\
        );

    \I__4098\ : InMux
    port map (
            O => \N__18574\,
            I => \N__18551\
        );

    \I__4097\ : Span4Mux_v
    port map (
            O => \N__18571\,
            I => \N__18546\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__18566\,
            I => \N__18546\
        );

    \I__4095\ : Span4Mux_h
    port map (
            O => \N__18561\,
            I => \N__18543\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__18558\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__18551\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__18546\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__18543\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__4090\ : InMux
    port map (
            O => \N__18534\,
            I => \N__18526\
        );

    \I__4089\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18526\
        );

    \I__4088\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18521\
        );

    \I__4087\ : InMux
    port map (
            O => \N__18531\,
            I => \N__18521\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__18526\,
            I => \N__18518\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__18521\,
            I => \N__18512\
        );

    \I__4084\ : Span4Mux_h
    port map (
            O => \N__18518\,
            I => \N__18509\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18517\,
            I => \N__18506\
        );

    \I__4082\ : InMux
    port map (
            O => \N__18516\,
            I => \N__18501\
        );

    \I__4081\ : InMux
    port map (
            O => \N__18515\,
            I => \N__18501\
        );

    \I__4080\ : Span4Mux_h
    port map (
            O => \N__18512\,
            I => \N__18496\
        );

    \I__4079\ : Span4Mux_h
    port map (
            O => \N__18509\,
            I => \N__18496\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__18506\,
            I => \Lab_UT.scdp.binValD_3\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__18501\,
            I => \Lab_UT.scdp.binValD_3\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__18496\,
            I => \Lab_UT.scdp.binValD_3\
        );

    \I__4075\ : InMux
    port map (
            O => \N__18489\,
            I => \N__18485\
        );

    \I__4074\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18479\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__18485\,
            I => \N__18476\
        );

    \I__4072\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18473\
        );

    \I__4071\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18468\
        );

    \I__4070\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18468\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__18479\,
            I => \Lab_UT.state_1_RNI2IGHH_0_0\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__18476\,
            I => \Lab_UT.state_1_RNI2IGHH_0_0\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__18473\,
            I => \Lab_UT.state_1_RNI2IGHH_0_0\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__18468\,
            I => \Lab_UT.state_1_RNI2IGHH_0_0\
        );

    \I__4065\ : InMux
    port map (
            O => \N__18459\,
            I => \N__18455\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__18458\,
            I => \N__18452\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__18455\,
            I => \N__18449\
        );

    \I__4062\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18446\
        );

    \I__4061\ : Odrv12
    port map (
            O => \N__18449\,
            I => \Lab_UT.scdp.key2_7\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__18446\,
            I => \Lab_UT.scdp.key2_7\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__18441\,
            I => \N__18434\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__18440\,
            I => \N__18424\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__18439\,
            I => \N__18421\
        );

    \I__4056\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18417\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18413\
        );

    \I__4054\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18410\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__18433\,
            I => \N__18407\
        );

    \I__4052\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18399\
        );

    \I__4051\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18399\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18430\,
            I => \N__18399\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__18429\,
            I => \N__18396\
        );

    \I__4048\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18392\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18387\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18387\
        );

    \I__4045\ : InMux
    port map (
            O => \N__18421\,
            I => \N__18382\
        );

    \I__4044\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18382\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__18417\,
            I => \N__18379\
        );

    \I__4042\ : InMux
    port map (
            O => \N__18416\,
            I => \N__18376\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__18413\,
            I => \N__18371\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__18410\,
            I => \N__18371\
        );

    \I__4039\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18366\
        );

    \I__4038\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18366\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__18399\,
            I => \N__18363\
        );

    \I__4036\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18360\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__18395\,
            I => \N__18357\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__18392\,
            I => \N__18352\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__18387\,
            I => \N__18347\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__18382\,
            I => \N__18347\
        );

    \I__4031\ : Span4Mux_s3_v
    port map (
            O => \N__18379\,
            I => \N__18338\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__18376\,
            I => \N__18338\
        );

    \I__4029\ : Span4Mux_h
    port map (
            O => \N__18371\,
            I => \N__18338\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__18366\,
            I => \N__18338\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__18363\,
            I => \N__18333\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__18360\,
            I => \N__18333\
        );

    \I__4025\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18330\
        );

    \I__4024\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18327\
        );

    \I__4023\ : CascadeMux
    port map (
            O => \N__18355\,
            I => \N__18324\
        );

    \I__4022\ : Span4Mux_v
    port map (
            O => \N__18352\,
            I => \N__18321\
        );

    \I__4021\ : Span4Mux_v
    port map (
            O => \N__18347\,
            I => \N__18318\
        );

    \I__4020\ : Span4Mux_v
    port map (
            O => \N__18338\,
            I => \N__18315\
        );

    \I__4019\ : Span4Mux_v
    port map (
            O => \N__18333\,
            I => \N__18312\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__18330\,
            I => \N__18307\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__18327\,
            I => \N__18307\
        );

    \I__4016\ : InMux
    port map (
            O => \N__18324\,
            I => \N__18304\
        );

    \I__4015\ : Sp12to4
    port map (
            O => \N__18321\,
            I => \N__18301\
        );

    \I__4014\ : Span4Mux_v
    port map (
            O => \N__18318\,
            I => \N__18296\
        );

    \I__4013\ : Span4Mux_s3_h
    port map (
            O => \N__18315\,
            I => \N__18296\
        );

    \I__4012\ : Span4Mux_s2_h
    port map (
            O => \N__18312\,
            I => \N__18291\
        );

    \I__4011\ : Span4Mux_v
    port map (
            O => \N__18307\,
            I => \N__18291\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__18304\,
            I => \Lab_UT.scctrl.state_i_1_0\
        );

    \I__4009\ : Odrv12
    port map (
            O => \N__18301\,
            I => \Lab_UT.scctrl.state_i_1_0\
        );

    \I__4008\ : Odrv4
    port map (
            O => \N__18296\,
            I => \Lab_UT.scctrl.state_i_1_0\
        );

    \I__4007\ : Odrv4
    port map (
            O => \N__18291\,
            I => \Lab_UT.scctrl.state_i_1_0\
        );

    \I__4006\ : InMux
    port map (
            O => \N__18282\,
            I => \N__18279\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__18279\,
            I => \N__18272\
        );

    \I__4004\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18269\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__18277\,
            I => \N__18266\
        );

    \I__4002\ : InMux
    port map (
            O => \N__18276\,
            I => \N__18260\
        );

    \I__4001\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18256\
        );

    \I__4000\ : Span4Mux_h
    port map (
            O => \N__18272\,
            I => \N__18251\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__18269\,
            I => \N__18251\
        );

    \I__3998\ : InMux
    port map (
            O => \N__18266\,
            I => \N__18248\
        );

    \I__3997\ : InMux
    port map (
            O => \N__18265\,
            I => \N__18242\
        );

    \I__3996\ : InMux
    port map (
            O => \N__18264\,
            I => \N__18239\
        );

    \I__3995\ : InMux
    port map (
            O => \N__18263\,
            I => \N__18235\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__18260\,
            I => \N__18232\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__18259\,
            I => \N__18227\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__18256\,
            I => \N__18222\
        );

    \I__3991\ : Span4Mux_v
    port map (
            O => \N__18251\,
            I => \N__18217\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__18248\,
            I => \N__18217\
        );

    \I__3989\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18212\
        );

    \I__3988\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18212\
        );

    \I__3987\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18209\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__18242\,
            I => \N__18204\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__18239\,
            I => \N__18204\
        );

    \I__3984\ : InMux
    port map (
            O => \N__18238\,
            I => \N__18200\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__18235\,
            I => \N__18197\
        );

    \I__3982\ : Span4Mux_s2_h
    port map (
            O => \N__18232\,
            I => \N__18194\
        );

    \I__3981\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18191\
        );

    \I__3980\ : InMux
    port map (
            O => \N__18230\,
            I => \N__18182\
        );

    \I__3979\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18182\
        );

    \I__3978\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18182\
        );

    \I__3977\ : InMux
    port map (
            O => \N__18225\,
            I => \N__18182\
        );

    \I__3976\ : Span4Mux_h
    port map (
            O => \N__18222\,
            I => \N__18177\
        );

    \I__3975\ : Span4Mux_h
    port map (
            O => \N__18217\,
            I => \N__18177\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__18212\,
            I => \N__18174\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__18209\,
            I => \N__18169\
        );

    \I__3972\ : Span12Mux_v
    port map (
            O => \N__18204\,
            I => \N__18169\
        );

    \I__3971\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18166\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__18200\,
            I => \Lab_UT.scctrl.N_296_i_0\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__18197\,
            I => \Lab_UT.scctrl.N_296_i_0\
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__18194\,
            I => \Lab_UT.scctrl.N_296_i_0\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__18191\,
            I => \Lab_UT.scctrl.N_296_i_0\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__18182\,
            I => \Lab_UT.scctrl.N_296_i_0\
        );

    \I__3965\ : Odrv4
    port map (
            O => \N__18177\,
            I => \Lab_UT.scctrl.N_296_i_0\
        );

    \I__3964\ : Odrv12
    port map (
            O => \N__18174\,
            I => \Lab_UT.scctrl.N_296_i_0\
        );

    \I__3963\ : Odrv12
    port map (
            O => \N__18169\,
            I => \Lab_UT.scctrl.N_296_i_0\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__18166\,
            I => \Lab_UT.scctrl.N_296_i_0\
        );

    \I__3961\ : InMux
    port map (
            O => \N__18147\,
            I => \N__18144\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__18144\,
            I => \N__18141\
        );

    \I__3959\ : Span4Mux_v
    port map (
            O => \N__18141\,
            I => \N__18138\
        );

    \I__3958\ : Span4Mux_h
    port map (
            O => \N__18138\,
            I => \N__18135\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__18135\,
            I => \Lab_UT.scctrl.next_state_RNO_1Z0Z_1\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__18132\,
            I => \Lab_UT.scctrl.N_319_cascade_\
        );

    \I__3955\ : InMux
    port map (
            O => \N__18129\,
            I => \N__18126\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__18126\,
            I => \N__18123\
        );

    \I__3953\ : Span4Mux_v
    port map (
            O => \N__18123\,
            I => \N__18120\
        );

    \I__3952\ : Odrv4
    port map (
            O => \N__18120\,
            I => \Lab_UT.scctrl.next_state_rst_1_0\
        );

    \I__3951\ : CascadeMux
    port map (
            O => \N__18117\,
            I => \Lab_UT.scctrl.N_414_cascade_\
        );

    \I__3950\ : InMux
    port map (
            O => \N__18114\,
            I => \N__18108\
        );

    \I__3949\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18108\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__18108\,
            I => \N__18105\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__18105\,
            I => \N__18102\
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__18102\,
            I => \Lab_UT.scctrl.next_state_rst_1_2\
        );

    \I__3945\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18096\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__18096\,
            I => \N__18093\
        );

    \I__3943\ : Span4Mux_h
    port map (
            O => \N__18093\,
            I => \N__18090\
        );

    \I__3942\ : Odrv4
    port map (
            O => \N__18090\,
            I => \Lab_UT.scctrl.N_319_1\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__18087\,
            I => \N__18082\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__18086\,
            I => \N__18079\
        );

    \I__3939\ : CascadeMux
    port map (
            O => \N__18085\,
            I => \N__18076\
        );

    \I__3938\ : InMux
    port map (
            O => \N__18082\,
            I => \N__18073\
        );

    \I__3937\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18068\
        );

    \I__3936\ : InMux
    port map (
            O => \N__18076\,
            I => \N__18062\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__18073\,
            I => \N__18059\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18072\,
            I => \N__18055\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__18071\,
            I => \N__18051\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__18068\,
            I => \N__18048\
        );

    \I__3931\ : InMux
    port map (
            O => \N__18067\,
            I => \N__18043\
        );

    \I__3930\ : InMux
    port map (
            O => \N__18066\,
            I => \N__18043\
        );

    \I__3929\ : InMux
    port map (
            O => \N__18065\,
            I => \N__18040\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__18062\,
            I => \N__18035\
        );

    \I__3927\ : Span4Mux_v
    port map (
            O => \N__18059\,
            I => \N__18032\
        );

    \I__3926\ : CascadeMux
    port map (
            O => \N__18058\,
            I => \N__18029\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__18055\,
            I => \N__18025\
        );

    \I__3924\ : CascadeMux
    port map (
            O => \N__18054\,
            I => \N__18022\
        );

    \I__3923\ : InMux
    port map (
            O => \N__18051\,
            I => \N__18019\
        );

    \I__3922\ : Span4Mux_h
    port map (
            O => \N__18048\,
            I => \N__18014\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__18043\,
            I => \N__18014\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__18040\,
            I => \N__18011\
        );

    \I__3919\ : InMux
    port map (
            O => \N__18039\,
            I => \N__18008\
        );

    \I__3918\ : InMux
    port map (
            O => \N__18038\,
            I => \N__18005\
        );

    \I__3917\ : Span4Mux_v
    port map (
            O => \N__18035\,
            I => \N__17999\
        );

    \I__3916\ : Span4Mux_s3_h
    port map (
            O => \N__18032\,
            I => \N__17999\
        );

    \I__3915\ : InMux
    port map (
            O => \N__18029\,
            I => \N__17994\
        );

    \I__3914\ : InMux
    port map (
            O => \N__18028\,
            I => \N__17994\
        );

    \I__3913\ : Span4Mux_s2_h
    port map (
            O => \N__18025\,
            I => \N__17991\
        );

    \I__3912\ : InMux
    port map (
            O => \N__18022\,
            I => \N__17988\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__18019\,
            I => \N__17983\
        );

    \I__3910\ : Span4Mux_s3_h
    port map (
            O => \N__18014\,
            I => \N__17983\
        );

    \I__3909\ : Span4Mux_v
    port map (
            O => \N__18011\,
            I => \N__17976\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__18008\,
            I => \N__17976\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__18005\,
            I => \N__17976\
        );

    \I__3906\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17973\
        );

    \I__3905\ : Span4Mux_v
    port map (
            O => \N__17999\,
            I => \N__17968\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__17994\,
            I => \N__17968\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__17991\,
            I => \Lab_UT.scctrl.state_2_rep2\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__17988\,
            I => \Lab_UT.scctrl.state_2_rep2\
        );

    \I__3901\ : Odrv4
    port map (
            O => \N__17983\,
            I => \Lab_UT.scctrl.state_2_rep2\
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__17976\,
            I => \Lab_UT.scctrl.state_2_rep2\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__17973\,
            I => \Lab_UT.scctrl.state_2_rep2\
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__17968\,
            I => \Lab_UT.scctrl.state_2_rep2\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__17955\,
            I => \Lab_UT.scctrl.N_7_1_cascade_\
        );

    \I__3896\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17945\
        );

    \I__3895\ : InMux
    port map (
            O => \N__17951\,
            I => \N__17936\
        );

    \I__3894\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17936\
        );

    \I__3893\ : InMux
    port map (
            O => \N__17949\,
            I => \N__17936\
        );

    \I__3892\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17936\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__17945\,
            I => \Lab_UT.state_ret_12_RNIUVHQG_0\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__17936\,
            I => \Lab_UT.state_ret_12_RNIUVHQG_0\
        );

    \I__3889\ : InMux
    port map (
            O => \N__17931\,
            I => \N__17927\
        );

    \I__3888\ : CascadeMux
    port map (
            O => \N__17930\,
            I => \N__17924\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__17927\,
            I => \N__17921\
        );

    \I__3886\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17918\
        );

    \I__3885\ : Odrv12
    port map (
            O => \N__17921\,
            I => \Lab_UT.scdp.key3_3\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__17918\,
            I => \Lab_UT.scdp.key3_3\
        );

    \I__3883\ : CascadeMux
    port map (
            O => \N__17913\,
            I => \N__17910\
        );

    \I__3882\ : InMux
    port map (
            O => \N__17910\,
            I => \N__17906\
        );

    \I__3881\ : InMux
    port map (
            O => \N__17909\,
            I => \N__17903\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__17906\,
            I => \Lab_UT.scdp.val_0_tz_3\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__17903\,
            I => \Lab_UT.scdp.val_0_tz_3\
        );

    \I__3878\ : CascadeMux
    port map (
            O => \N__17898\,
            I => \N__17887\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__17897\,
            I => \N__17881\
        );

    \I__3876\ : CascadeMux
    port map (
            O => \N__17896\,
            I => \N__17878\
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__17895\,
            I => \N__17875\
        );

    \I__3874\ : CascadeMux
    port map (
            O => \N__17894\,
            I => \N__17872\
        );

    \I__3873\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17869\
        );

    \I__3872\ : InMux
    port map (
            O => \N__17892\,
            I => \N__17866\
        );

    \I__3871\ : InMux
    port map (
            O => \N__17891\,
            I => \N__17859\
        );

    \I__3870\ : InMux
    port map (
            O => \N__17890\,
            I => \N__17859\
        );

    \I__3869\ : InMux
    port map (
            O => \N__17887\,
            I => \N__17859\
        );

    \I__3868\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17856\
        );

    \I__3867\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17852\
        );

    \I__3866\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17841\
        );

    \I__3865\ : InMux
    port map (
            O => \N__17881\,
            I => \N__17841\
        );

    \I__3864\ : InMux
    port map (
            O => \N__17878\,
            I => \N__17841\
        );

    \I__3863\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17841\
        );

    \I__3862\ : InMux
    port map (
            O => \N__17872\,
            I => \N__17841\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__17869\,
            I => \N__17834\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__17866\,
            I => \N__17834\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__17859\,
            I => \N__17834\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__17856\,
            I => \N__17831\
        );

    \I__3857\ : InMux
    port map (
            O => \N__17855\,
            I => \N__17828\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__17852\,
            I => \N__17820\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__17841\,
            I => \N__17820\
        );

    \I__3854\ : Span4Mux_h
    port map (
            O => \N__17834\,
            I => \N__17820\
        );

    \I__3853\ : Span4Mux_h
    port map (
            O => \N__17831\,
            I => \N__17817\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__17828\,
            I => \N__17814\
        );

    \I__3851\ : InMux
    port map (
            O => \N__17827\,
            I => \N__17811\
        );

    \I__3850\ : Span4Mux_v
    port map (
            O => \N__17820\,
            I => \N__17808\
        );

    \I__3849\ : Span4Mux_v
    port map (
            O => \N__17817\,
            I => \N__17801\
        );

    \I__3848\ : Span4Mux_h
    port map (
            O => \N__17814\,
            I => \N__17801\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__17811\,
            I => \N__17801\
        );

    \I__3846\ : Span4Mux_h
    port map (
            O => \N__17808\,
            I => \N__17798\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__17801\,
            I => bu_rx_data_i_2_3
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__17798\,
            I => bu_rx_data_i_2_3
        );

    \I__3843\ : InMux
    port map (
            O => \N__17793\,
            I => \N__17788\
        );

    \I__3842\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17785\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__17791\,
            I => \N__17782\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__17788\,
            I => \N__17779\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__17785\,
            I => \N__17776\
        );

    \I__3838\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17773\
        );

    \I__3837\ : Span4Mux_h
    port map (
            O => \N__17779\,
            I => \N__17768\
        );

    \I__3836\ : Span4Mux_v
    port map (
            O => \N__17776\,
            I => \N__17768\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__17773\,
            I => \buart.Z_rx.N_301\
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__17768\,
            I => \buart.Z_rx.N_301\
        );

    \I__3833\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17759\
        );

    \I__3832\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17756\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__17759\,
            I => \N__17753\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__17756\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__3829\ : Odrv12
    port map (
            O => \N__17753\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__17748\,
            I => \N__17744\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17736\
        );

    \I__3826\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17736\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17743\,
            I => \N__17736\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__17736\,
            I => \N__17731\
        );

    \I__3823\ : InMux
    port map (
            O => \N__17735\,
            I => \N__17728\
        );

    \I__3822\ : InMux
    port map (
            O => \N__17734\,
            I => \N__17725\
        );

    \I__3821\ : Span4Mux_v
    port map (
            O => \N__17731\,
            I => \N__17720\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__17728\,
            I => \N__17720\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__17725\,
            I => \N__17717\
        );

    \I__3818\ : Span4Mux_h
    port map (
            O => \N__17720\,
            I => \N__17714\
        );

    \I__3817\ : Span4Mux_h
    port map (
            O => \N__17717\,
            I => \N__17711\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__17714\,
            I => \N__17708\
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__17711\,
            I => \buart__rx_hh_1\
        );

    \I__3814\ : Odrv4
    port map (
            O => \N__17708\,
            I => \buart__rx_hh_1\
        );

    \I__3813\ : InMux
    port map (
            O => \N__17703\,
            I => \N__17691\
        );

    \I__3812\ : InMux
    port map (
            O => \N__17702\,
            I => \N__17686\
        );

    \I__3811\ : InMux
    port map (
            O => \N__17701\,
            I => \N__17686\
        );

    \I__3810\ : CascadeMux
    port map (
            O => \N__17700\,
            I => \N__17682\
        );

    \I__3809\ : CascadeMux
    port map (
            O => \N__17699\,
            I => \N__17679\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__17698\,
            I => \N__17676\
        );

    \I__3807\ : InMux
    port map (
            O => \N__17697\,
            I => \N__17666\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17696\,
            I => \N__17666\
        );

    \I__3805\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17666\
        );

    \I__3804\ : InMux
    port map (
            O => \N__17694\,
            I => \N__17666\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__17691\,
            I => \N__17661\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__17686\,
            I => \N__17661\
        );

    \I__3801\ : InMux
    port map (
            O => \N__17685\,
            I => \N__17652\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17682\,
            I => \N__17652\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17679\,
            I => \N__17652\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17676\,
            I => \N__17652\
        );

    \I__3797\ : InMux
    port map (
            O => \N__17675\,
            I => \N__17649\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__17666\,
            I => \N__17646\
        );

    \I__3795\ : Span4Mux_v
    port map (
            O => \N__17661\,
            I => \N__17641\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__17652\,
            I => \N__17641\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__17649\,
            I => \N__17634\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__17646\,
            I => \N__17634\
        );

    \I__3791\ : Span4Mux_h
    port map (
            O => \N__17641\,
            I => \N__17634\
        );

    \I__3790\ : Span4Mux_h
    port map (
            O => \N__17634\,
            I => \N__17631\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__17631\,
            I => \buart.Z_rx.startbit\
        );

    \I__3788\ : InMux
    port map (
            O => \N__17628\,
            I => \N__17623\
        );

    \I__3787\ : InMux
    port map (
            O => \N__17627\,
            I => \N__17618\
        );

    \I__3786\ : InMux
    port map (
            O => \N__17626\,
            I => \N__17618\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17623\,
            I => \N__17610\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__17618\,
            I => \N__17610\
        );

    \I__3783\ : InMux
    port map (
            O => \N__17617\,
            I => \N__17605\
        );

    \I__3782\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17605\
        );

    \I__3781\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17602\
        );

    \I__3780\ : Span4Mux_v
    port map (
            O => \N__17610\,
            I => \N__17597\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__17605\,
            I => \N__17594\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__17602\,
            I => \N__17591\
        );

    \I__3777\ : InMux
    port map (
            O => \N__17601\,
            I => \N__17586\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17600\,
            I => \N__17586\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__17597\,
            I => \Lab_UT.scdp.binValD_0\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__17594\,
            I => \Lab_UT.scdp.binValD_0\
        );

    \I__3773\ : Odrv4
    port map (
            O => \N__17591\,
            I => \Lab_UT.scdp.binValD_0\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__17586\,
            I => \Lab_UT.scdp.binValD_0\
        );

    \I__3771\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17574\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__17574\,
            I => \N__17570\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__17573\,
            I => \N__17567\
        );

    \I__3768\ : Span4Mux_v
    port map (
            O => \N__17570\,
            I => \N__17564\
        );

    \I__3767\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17561\
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__17564\,
            I => \Lab_UT.scdp.key0_0\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__17561\,
            I => \Lab_UT.scdp.key0_0\
        );

    \I__3764\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17550\
        );

    \I__3763\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17550\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__17550\,
            I => \N__17546\
        );

    \I__3761\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17541\
        );

    \I__3760\ : Span4Mux_h
    port map (
            O => \N__17546\,
            I => \N__17538\
        );

    \I__3759\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17533\
        );

    \I__3758\ : InMux
    port map (
            O => \N__17544\,
            I => \N__17533\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__17541\,
            I => \Lab_UT.state_1_RNIO1RJH_0_2\
        );

    \I__3756\ : Odrv4
    port map (
            O => \N__17538\,
            I => \Lab_UT.state_1_RNIO1RJH_0_2\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__17533\,
            I => \Lab_UT.state_1_RNIO1RJH_0_2\
        );

    \I__3754\ : InMux
    port map (
            O => \N__17526\,
            I => \N__17522\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__17525\,
            I => \N__17519\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__17522\,
            I => \N__17516\
        );

    \I__3751\ : InMux
    port map (
            O => \N__17519\,
            I => \N__17513\
        );

    \I__3750\ : Odrv12
    port map (
            O => \N__17516\,
            I => \Lab_UT.scdp.key0_1\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__17513\,
            I => \Lab_UT.scdp.key0_1\
        );

    \I__3748\ : InMux
    port map (
            O => \N__17508\,
            I => \N__17501\
        );

    \I__3747\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17498\
        );

    \I__3746\ : InMux
    port map (
            O => \N__17506\,
            I => \N__17493\
        );

    \I__3745\ : InMux
    port map (
            O => \N__17505\,
            I => \N__17493\
        );

    \I__3744\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17490\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__17501\,
            I => \Lab_UT.state_1_ret_3_RNI23U7H_0\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__17498\,
            I => \Lab_UT.state_1_ret_3_RNI23U7H_0\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__17493\,
            I => \Lab_UT.state_1_ret_3_RNI23U7H_0\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__17490\,
            I => \Lab_UT.state_1_ret_3_RNI23U7H_0\
        );

    \I__3739\ : InMux
    port map (
            O => \N__17481\,
            I => \N__17478\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__17478\,
            I => \N__17475\
        );

    \I__3737\ : Span4Mux_v
    port map (
            O => \N__17475\,
            I => \N__17471\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__17474\,
            I => \N__17468\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__17471\,
            I => \N__17465\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17468\,
            I => \N__17462\
        );

    \I__3733\ : Odrv4
    port map (
            O => \N__17465\,
            I => \Lab_UT.scdp.key1_5\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__17462\,
            I => \Lab_UT.scdp.key1_5\
        );

    \I__3731\ : InMux
    port map (
            O => \N__17457\,
            I => \N__17450\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17456\,
            I => \N__17447\
        );

    \I__3729\ : InMux
    port map (
            O => \N__17455\,
            I => \N__17444\
        );

    \I__3728\ : InMux
    port map (
            O => \N__17454\,
            I => \N__17439\
        );

    \I__3727\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17439\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__17450\,
            I => \Lab_UT.state_ret_RNIK5UKH_0\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__17447\,
            I => \Lab_UT.state_ret_RNIK5UKH_0\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__17444\,
            I => \Lab_UT.state_ret_RNIK5UKH_0\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__17439\,
            I => \Lab_UT.state_ret_RNIK5UKH_0\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17430\,
            I => \N__17427\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__17427\,
            I => \N__17423\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__17426\,
            I => \N__17420\
        );

    \I__3719\ : Span4Mux_h
    port map (
            O => \N__17423\,
            I => \N__17417\
        );

    \I__3718\ : InMux
    port map (
            O => \N__17420\,
            I => \N__17414\
        );

    \I__3717\ : Odrv4
    port map (
            O => \N__17417\,
            I => \Lab_UT.scdp.key2_3\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__17414\,
            I => \Lab_UT.scdp.key2_3\
        );

    \I__3715\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17403\
        );

    \I__3714\ : InMux
    port map (
            O => \N__17408\,
            I => \N__17403\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__17403\,
            I => \N__17399\
        );

    \I__3712\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17396\
        );

    \I__3711\ : Span4Mux_v
    port map (
            O => \N__17399\,
            I => \N__17388\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__17396\,
            I => \N__17388\
        );

    \I__3709\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17381\
        );

    \I__3708\ : InMux
    port map (
            O => \N__17394\,
            I => \N__17381\
        );

    \I__3707\ : InMux
    port map (
            O => \N__17393\,
            I => \N__17381\
        );

    \I__3706\ : Span4Mux_h
    port map (
            O => \N__17388\,
            I => \N__17376\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__17381\,
            I => \N__17376\
        );

    \I__3704\ : Span4Mux_v
    port map (
            O => \N__17376\,
            I => \N__17371\
        );

    \I__3703\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17366\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17366\
        );

    \I__3701\ : Span4Mux_s3_h
    port map (
            O => \N__17371\,
            I => \N__17363\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__17366\,
            I => \Lab_UT.scdp.binValD_1\
        );

    \I__3699\ : Odrv4
    port map (
            O => \N__17363\,
            I => \Lab_UT.scdp.binValD_1\
        );

    \I__3698\ : InMux
    port map (
            O => \N__17358\,
            I => \N__17351\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17357\,
            I => \N__17348\
        );

    \I__3696\ : InMux
    port map (
            O => \N__17356\,
            I => \N__17341\
        );

    \I__3695\ : InMux
    port map (
            O => \N__17355\,
            I => \N__17341\
        );

    \I__3694\ : InMux
    port map (
            O => \N__17354\,
            I => \N__17341\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__17351\,
            I => \Lab_UT.state_ret_12_RNI2SEPG_0\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__17348\,
            I => \Lab_UT.state_ret_12_RNI2SEPG_0\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__17341\,
            I => \Lab_UT.state_ret_12_RNI2SEPG_0\
        );

    \I__3690\ : InMux
    port map (
            O => \N__17334\,
            I => \N__17331\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__17331\,
            I => \N__17327\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__17330\,
            I => \N__17324\
        );

    \I__3687\ : Span4Mux_s2_v
    port map (
            O => \N__17327\,
            I => \N__17321\
        );

    \I__3686\ : InMux
    port map (
            O => \N__17324\,
            I => \N__17318\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__17321\,
            I => \Lab_UT.scdp.key1_1\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__17318\,
            I => \Lab_UT.scdp.key1_1\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__17313\,
            I => \Lab_UT.scdp.N_378_cascade_\
        );

    \I__3682\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17307\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__17307\,
            I => \N__17303\
        );

    \I__3680\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17300\
        );

    \I__3679\ : Span4Mux_h
    port map (
            O => \N__17303\,
            I => \N__17297\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__17300\,
            I => \Lab_UT.scdp.byteToDecrypt_4\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__17297\,
            I => \Lab_UT.scdp.byteToDecrypt_4\
        );

    \I__3676\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17288\
        );

    \I__3675\ : InMux
    port map (
            O => \N__17291\,
            I => \N__17285\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__17288\,
            I => \Lab_UT.scdp.val_i_0_0\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__17285\,
            I => \Lab_UT.scdp.val_i_0_0\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__17280\,
            I => \N__17277\
        );

    \I__3671\ : InMux
    port map (
            O => \N__17277\,
            I => \N__17271\
        );

    \I__3670\ : InMux
    port map (
            O => \N__17276\,
            I => \N__17271\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__17271\,
            I => \Lab_UT.scdp.N_378\
        );

    \I__3668\ : CascadeMux
    port map (
            O => \N__17268\,
            I => \N__17264\
        );

    \I__3667\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17259\
        );

    \I__3666\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17252\
        );

    \I__3665\ : InMux
    port map (
            O => \N__17263\,
            I => \N__17252\
        );

    \I__3664\ : InMux
    port map (
            O => \N__17262\,
            I => \N__17252\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__17259\,
            I => \N__17248\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__17252\,
            I => \N__17245\
        );

    \I__3661\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17242\
        );

    \I__3660\ : Span4Mux_h
    port map (
            O => \N__17248\,
            I => \N__17237\
        );

    \I__3659\ : Span4Mux_v
    port map (
            O => \N__17245\,
            I => \N__17237\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__17242\,
            I => \Lab_UT.scdp.u1.byteToDecryptZ0Z_0\
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__17237\,
            I => \Lab_UT.scdp.u1.byteToDecryptZ0Z_0\
        );

    \I__3656\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17229\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__17229\,
            I => \N__17226\
        );

    \I__3654\ : Span4Mux_v
    port map (
            O => \N__17226\,
            I => \N__17223\
        );

    \I__3653\ : Span4Mux_h
    port map (
            O => \N__17223\,
            I => \N__17220\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__17220\,
            I => \Lab_UT.scdp.a2b.val_0_tz_0_3\
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__17217\,
            I => \N__17214\
        );

    \I__3650\ : InMux
    port map (
            O => \N__17214\,
            I => \N__17207\
        );

    \I__3649\ : InMux
    port map (
            O => \N__17213\,
            I => \N__17207\
        );

    \I__3648\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17202\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__17207\,
            I => \N__17199\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__17206\,
            I => \N__17192\
        );

    \I__3645\ : InMux
    port map (
            O => \N__17205\,
            I => \N__17187\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__17202\,
            I => \N__17182\
        );

    \I__3643\ : Span4Mux_s3_v
    port map (
            O => \N__17199\,
            I => \N__17182\
        );

    \I__3642\ : InMux
    port map (
            O => \N__17198\,
            I => \N__17175\
        );

    \I__3641\ : InMux
    port map (
            O => \N__17197\,
            I => \N__17175\
        );

    \I__3640\ : InMux
    port map (
            O => \N__17196\,
            I => \N__17175\
        );

    \I__3639\ : InMux
    port map (
            O => \N__17195\,
            I => \N__17172\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17167\
        );

    \I__3637\ : InMux
    port map (
            O => \N__17191\,
            I => \N__17167\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__17190\,
            I => \N__17156\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__17187\,
            I => \N__17152\
        );

    \I__3634\ : Span4Mux_v
    port map (
            O => \N__17182\,
            I => \N__17147\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__17175\,
            I => \N__17147\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__17172\,
            I => \N__17142\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__17167\,
            I => \N__17142\
        );

    \I__3630\ : InMux
    port map (
            O => \N__17166\,
            I => \N__17133\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17165\,
            I => \N__17133\
        );

    \I__3628\ : InMux
    port map (
            O => \N__17164\,
            I => \N__17133\
        );

    \I__3627\ : InMux
    port map (
            O => \N__17163\,
            I => \N__17133\
        );

    \I__3626\ : InMux
    port map (
            O => \N__17162\,
            I => \N__17130\
        );

    \I__3625\ : InMux
    port map (
            O => \N__17161\,
            I => \N__17125\
        );

    \I__3624\ : InMux
    port map (
            O => \N__17160\,
            I => \N__17118\
        );

    \I__3623\ : InMux
    port map (
            O => \N__17159\,
            I => \N__17118\
        );

    \I__3622\ : InMux
    port map (
            O => \N__17156\,
            I => \N__17118\
        );

    \I__3621\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17115\
        );

    \I__3620\ : Span4Mux_v
    port map (
            O => \N__17152\,
            I => \N__17110\
        );

    \I__3619\ : Span4Mux_v
    port map (
            O => \N__17147\,
            I => \N__17110\
        );

    \I__3618\ : Span4Mux_v
    port map (
            O => \N__17142\,
            I => \N__17107\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__17133\,
            I => \N__17102\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__17130\,
            I => \N__17102\
        );

    \I__3615\ : InMux
    port map (
            O => \N__17129\,
            I => \N__17099\
        );

    \I__3614\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17096\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__17125\,
            I => \N__17091\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__17118\,
            I => \N__17091\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__17115\,
            I => bu_rx_data_1
        );

    \I__3610\ : Odrv4
    port map (
            O => \N__17110\,
            I => bu_rx_data_1
        );

    \I__3609\ : Odrv4
    port map (
            O => \N__17107\,
            I => bu_rx_data_1
        );

    \I__3608\ : Odrv12
    port map (
            O => \N__17102\,
            I => bu_rx_data_1
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__17099\,
            I => bu_rx_data_1
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__17096\,
            I => bu_rx_data_1
        );

    \I__3605\ : Odrv4
    port map (
            O => \N__17091\,
            I => bu_rx_data_1
        );

    \I__3604\ : CascadeMux
    port map (
            O => \N__17076\,
            I => \N__17071\
        );

    \I__3603\ : InMux
    port map (
            O => \N__17075\,
            I => \N__17064\
        );

    \I__3602\ : InMux
    port map (
            O => \N__17074\,
            I => \N__17064\
        );

    \I__3601\ : InMux
    port map (
            O => \N__17071\,
            I => \N__17064\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__17064\,
            I => \N__17061\
        );

    \I__3599\ : Span4Mux_v
    port map (
            O => \N__17061\,
            I => \N__17058\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__17058\,
            I => bu_rx_data_i_2_2
        );

    \I__3597\ : InMux
    port map (
            O => \N__17055\,
            I => \N__17044\
        );

    \I__3596\ : InMux
    port map (
            O => \N__17054\,
            I => \N__17044\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__17053\,
            I => \N__17038\
        );

    \I__3594\ : InMux
    port map (
            O => \N__17052\,
            I => \N__17027\
        );

    \I__3593\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17027\
        );

    \I__3592\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17027\
        );

    \I__3591\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17027\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__17044\,
            I => \N__17024\
        );

    \I__3589\ : InMux
    port map (
            O => \N__17043\,
            I => \N__17019\
        );

    \I__3588\ : InMux
    port map (
            O => \N__17042\,
            I => \N__17008\
        );

    \I__3587\ : InMux
    port map (
            O => \N__17041\,
            I => \N__17008\
        );

    \I__3586\ : InMux
    port map (
            O => \N__17038\,
            I => \N__17008\
        );

    \I__3585\ : InMux
    port map (
            O => \N__17037\,
            I => \N__17008\
        );

    \I__3584\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17008\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__17027\,
            I => \N__17005\
        );

    \I__3582\ : Span4Mux_v
    port map (
            O => \N__17024\,
            I => \N__17002\
        );

    \I__3581\ : InMux
    port map (
            O => \N__17023\,
            I => \N__16997\
        );

    \I__3580\ : InMux
    port map (
            O => \N__17022\,
            I => \N__16997\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__17019\,
            I => \N__16992\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__17008\,
            I => \N__16992\
        );

    \I__3577\ : Span4Mux_v
    port map (
            O => \N__17005\,
            I => \N__16983\
        );

    \I__3576\ : Span4Mux_h
    port map (
            O => \N__17002\,
            I => \N__16983\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__16997\,
            I => \N__16980\
        );

    \I__3574\ : Span4Mux_v
    port map (
            O => \N__16992\,
            I => \N__16977\
        );

    \I__3573\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16972\
        );

    \I__3572\ : InMux
    port map (
            O => \N__16990\,
            I => \N__16972\
        );

    \I__3571\ : InMux
    port map (
            O => \N__16989\,
            I => \N__16967\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16988\,
            I => \N__16967\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__16983\,
            I => bu_rx_data_i_2_0
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__16980\,
            I => bu_rx_data_i_2_0
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__16977\,
            I => bu_rx_data_i_2_0
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__16972\,
            I => bu_rx_data_i_2_0
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__16967\,
            I => bu_rx_data_i_2_0
        );

    \I__3564\ : InMux
    port map (
            O => \N__16956\,
            I => \N__16953\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__16953\,
            I => \N__16948\
        );

    \I__3562\ : InMux
    port map (
            O => \N__16952\,
            I => \N__16943\
        );

    \I__3561\ : InMux
    port map (
            O => \N__16951\,
            I => \N__16943\
        );

    \I__3560\ : Span4Mux_v
    port map (
            O => \N__16948\,
            I => \N__16940\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__16943\,
            I => \N__16937\
        );

    \I__3558\ : Odrv4
    port map (
            O => \N__16940\,
            I => \Lab_UT.sccDnibble1En\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__16937\,
            I => \Lab_UT.sccDnibble1En\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__16932\,
            I => \Lab_UT.scdp.val_0_tz_3_cascade_\
        );

    \I__3555\ : InMux
    port map (
            O => \N__16929\,
            I => \N__16919\
        );

    \I__3554\ : InMux
    port map (
            O => \N__16928\,
            I => \N__16919\
        );

    \I__3553\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16919\
        );

    \I__3552\ : InMux
    port map (
            O => \N__16926\,
            I => \N__16916\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__16919\,
            I => \N__16913\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__16916\,
            I => \Lab_UT.scdp.byteToDecrypt_7\
        );

    \I__3549\ : Odrv12
    port map (
            O => \N__16913\,
            I => \Lab_UT.scdp.byteToDecrypt_7\
        );

    \I__3548\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16904\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__16907\,
            I => \N__16901\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__16904\,
            I => \N__16898\
        );

    \I__3545\ : InMux
    port map (
            O => \N__16901\,
            I => \N__16895\
        );

    \I__3544\ : Odrv12
    port map (
            O => \N__16898\,
            I => \Lab_UT.scdp.key2_0\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__16895\,
            I => \Lab_UT.scdp.key2_0\
        );

    \I__3542\ : InMux
    port map (
            O => \N__16890\,
            I => \N__16887\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__16887\,
            I => \N__16883\
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__16886\,
            I => \N__16880\
        );

    \I__3539\ : Span12Mux_s3_v
    port map (
            O => \N__16883\,
            I => \N__16877\
        );

    \I__3538\ : InMux
    port map (
            O => \N__16880\,
            I => \N__16874\
        );

    \I__3537\ : Odrv12
    port map (
            O => \N__16877\,
            I => \Lab_UT.scdp.key2_1\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__16874\,
            I => \Lab_UT.scdp.key2_1\
        );

    \I__3535\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16865\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__16868\,
            I => \N__16862\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__16865\,
            I => \N__16859\
        );

    \I__3532\ : InMux
    port map (
            O => \N__16862\,
            I => \N__16856\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__16859\,
            I => \Lab_UT.scdp.key3_0\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__16856\,
            I => \Lab_UT.scdp.key3_0\
        );

    \I__3529\ : InMux
    port map (
            O => \N__16851\,
            I => \N__16848\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__16848\,
            I => \N__16845\
        );

    \I__3527\ : Span4Mux_h
    port map (
            O => \N__16845\,
            I => \N__16841\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__16844\,
            I => \N__16838\
        );

    \I__3525\ : Span4Mux_h
    port map (
            O => \N__16841\,
            I => \N__16835\
        );

    \I__3524\ : InMux
    port map (
            O => \N__16838\,
            I => \N__16832\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__16835\,
            I => \Lab_UT.scdp.key3_1\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__16832\,
            I => \Lab_UT.scdp.key3_1\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__16827\,
            I => \N__16821\
        );

    \I__3520\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16817\
        );

    \I__3519\ : InMux
    port map (
            O => \N__16825\,
            I => \N__16808\
        );

    \I__3518\ : InMux
    port map (
            O => \N__16824\,
            I => \N__16808\
        );

    \I__3517\ : InMux
    port map (
            O => \N__16821\,
            I => \N__16808\
        );

    \I__3516\ : InMux
    port map (
            O => \N__16820\,
            I => \N__16808\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__16817\,
            I => \N__16805\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__16808\,
            I => \N__16802\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__16805\,
            I => \N__16796\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__16802\,
            I => \N__16793\
        );

    \I__3511\ : InMux
    port map (
            O => \N__16801\,
            I => \N__16790\
        );

    \I__3510\ : InMux
    port map (
            O => \N__16800\,
            I => \N__16785\
        );

    \I__3509\ : InMux
    port map (
            O => \N__16799\,
            I => \N__16785\
        );

    \I__3508\ : Odrv4
    port map (
            O => \N__16796\,
            I => \Lab_UT.scdp.binValD_2\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__16793\,
            I => \Lab_UT.scdp.binValD_2\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__16790\,
            I => \Lab_UT.scdp.binValD_2\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__16785\,
            I => \Lab_UT.scdp.binValD_2\
        );

    \I__3504\ : InMux
    port map (
            O => \N__16776\,
            I => \N__16773\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__16773\,
            I => \N__16769\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__16772\,
            I => \N__16766\
        );

    \I__3501\ : Span4Mux_s3_v
    port map (
            O => \N__16769\,
            I => \N__16763\
        );

    \I__3500\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16760\
        );

    \I__3499\ : Odrv4
    port map (
            O => \N__16763\,
            I => \Lab_UT.scdp.key3_2\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__16760\,
            I => \Lab_UT.scdp.key3_2\
        );

    \I__3497\ : InMux
    port map (
            O => \N__16755\,
            I => \N__16752\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__16752\,
            I => \N__16749\
        );

    \I__3495\ : Span4Mux_v
    port map (
            O => \N__16749\,
            I => \N__16746\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__16746\,
            I => \Lab_UT.scctrl.g1_1_0\
        );

    \I__3493\ : InMux
    port map (
            O => \N__16743\,
            I => \N__16740\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__16740\,
            I => \Lab_UT.scctrl.N_444_1_0\
        );

    \I__3491\ : InMux
    port map (
            O => \N__16737\,
            I => \N__16731\
        );

    \I__3490\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16731\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__16731\,
            I => \N__16727\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16730\,
            I => \N__16724\
        );

    \I__3487\ : Odrv4
    port map (
            O => \N__16727\,
            I => \Lab_UT.scctrl.g0_1_1\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__16724\,
            I => \Lab_UT.scctrl.g0_1_1\
        );

    \I__3485\ : CascadeMux
    port map (
            O => \N__16719\,
            I => \Lab_UT.scctrl.g1_0_3_cascade_\
        );

    \I__3484\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16713\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__16713\,
            I => \Lab_UT.scctrl.g1_2\
        );

    \I__3482\ : InMux
    port map (
            O => \N__16710\,
            I => \N__16707\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__16707\,
            I => \Lab_UT.scctrl.N_418_0_0\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__16704\,
            I => \N__16700\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16697\
        );

    \I__3478\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16694\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__16697\,
            I => \N__16691\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__16694\,
            I => \N__16688\
        );

    \I__3475\ : Span4Mux_v
    port map (
            O => \N__16691\,
            I => \N__16685\
        );

    \I__3474\ : Span4Mux_v
    port map (
            O => \N__16688\,
            I => \N__16682\
        );

    \I__3473\ : Odrv4
    port map (
            O => \N__16685\,
            I => \Lab_UT.scctrl.g0_0\
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__16682\,
            I => \Lab_UT.scctrl.g0_0\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16674\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__16674\,
            I => \Lab_UT.scctrl.g0_2_1\
        );

    \I__3469\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16668\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__16668\,
            I => \Lab_UT.scctrl.g0_9_a2_2\
        );

    \I__3467\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16662\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__16662\,
            I => \N__16658\
        );

    \I__3465\ : InMux
    port map (
            O => \N__16661\,
            I => \N__16655\
        );

    \I__3464\ : Span12Mux_s4_v
    port map (
            O => \N__16658\,
            I => \N__16652\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__16655\,
            I => \Lab_UT.scdp.byteToDecrypt_3\
        );

    \I__3462\ : Odrv12
    port map (
            O => \N__16652\,
            I => \Lab_UT.scdp.byteToDecrypt_3\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__16647\,
            I => \Lab_UT.scdp.val_i_0_0_cascade_\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16635\
        );

    \I__3459\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16632\
        );

    \I__3458\ : InMux
    port map (
            O => \N__16642\,
            I => \N__16629\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__16641\,
            I => \N__16626\
        );

    \I__3456\ : CascadeMux
    port map (
            O => \N__16640\,
            I => \N__16623\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__16639\,
            I => \N__16620\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__16638\,
            I => \N__16617\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__16635\,
            I => \N__16612\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__16632\,
            I => \N__16612\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__16629\,
            I => \N__16609\
        );

    \I__3450\ : InMux
    port map (
            O => \N__16626\,
            I => \N__16604\
        );

    \I__3449\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16604\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16620\,
            I => \N__16599\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16617\,
            I => \N__16599\
        );

    \I__3446\ : Span4Mux_v
    port map (
            O => \N__16612\,
            I => \N__16596\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__16609\,
            I => \N__16589\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__16604\,
            I => \N__16589\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__16599\,
            I => \N__16589\
        );

    \I__3442\ : Span4Mux_v
    port map (
            O => \N__16596\,
            I => \N__16584\
        );

    \I__3441\ : Span4Mux_v
    port map (
            O => \N__16589\,
            I => \N__16584\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__16584\,
            I => \Lab_UT.scdp.a2b.N_280\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__16581\,
            I => \N__16577\
        );

    \I__3438\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16572\
        );

    \I__3437\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16569\
        );

    \I__3436\ : InMux
    port map (
            O => \N__16576\,
            I => \N__16566\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__16575\,
            I => \N__16563\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__16572\,
            I => \N__16556\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__16569\,
            I => \N__16553\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__16566\,
            I => \N__16550\
        );

    \I__3431\ : InMux
    port map (
            O => \N__16563\,
            I => \N__16547\
        );

    \I__3430\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16544\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16561\,
            I => \N__16539\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16560\,
            I => \N__16539\
        );

    \I__3427\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16536\
        );

    \I__3426\ : Span4Mux_v
    port map (
            O => \N__16556\,
            I => \N__16533\
        );

    \I__3425\ : Span4Mux_v
    port map (
            O => \N__16553\,
            I => \N__16530\
        );

    \I__3424\ : Span4Mux_h
    port map (
            O => \N__16550\,
            I => \N__16527\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__16547\,
            I => \N__16524\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__16544\,
            I => \N__16521\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__16539\,
            I => \N__16516\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__16536\,
            I => \N__16516\
        );

    \I__3419\ : Span4Mux_h
    port map (
            O => \N__16533\,
            I => \N__16507\
        );

    \I__3418\ : Span4Mux_s2_h
    port map (
            O => \N__16530\,
            I => \N__16507\
        );

    \I__3417\ : Span4Mux_v
    port map (
            O => \N__16527\,
            I => \N__16507\
        );

    \I__3416\ : Span4Mux_v
    port map (
            O => \N__16524\,
            I => \N__16507\
        );

    \I__3415\ : Span4Mux_v
    port map (
            O => \N__16521\,
            I => \N__16502\
        );

    \I__3414\ : Span4Mux_v
    port map (
            O => \N__16516\,
            I => \N__16502\
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__16507\,
            I => bu_rx_data_0
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__16502\,
            I => bu_rx_data_0
        );

    \I__3411\ : CEMux
    port map (
            O => \N__16497\,
            I => \N__16494\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__16494\,
            I => \N__16491\
        );

    \I__3409\ : Span4Mux_v
    port map (
            O => \N__16491\,
            I => \N__16488\
        );

    \I__3408\ : Odrv4
    port map (
            O => \N__16488\,
            I => \Lab_UT.scctrl.N_398i_i\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__16485\,
            I => \N__16482\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16479\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__16479\,
            I => \N__16476\
        );

    \I__3404\ : Span4Mux_v
    port map (
            O => \N__16476\,
            I => \N__16473\
        );

    \I__3403\ : Span4Mux_h
    port map (
            O => \N__16473\,
            I => \N__16470\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__16470\,
            I => \Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0_0\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16461\
        );

    \I__3400\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16461\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__16461\,
            I => \Lab_UT.scctrl.nibbleInZ0Z1\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__16458\,
            I => \Lab_UT.scctrl.N_69_cascade_\
        );

    \I__3397\ : CascadeMux
    port map (
            O => \N__16455\,
            I => \Lab_UT.sccDnibble1En_cascade_\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16452\,
            I => \N__16448\
        );

    \I__3395\ : IoInMux
    port map (
            O => \N__16451\,
            I => \N__16444\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__16448\,
            I => \N__16441\
        );

    \I__3393\ : InMux
    port map (
            O => \N__16447\,
            I => \N__16438\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__16444\,
            I => \N__16435\
        );

    \I__3391\ : Span4Mux_h
    port map (
            O => \N__16441\,
            I => \N__16432\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__16438\,
            I => \N__16429\
        );

    \I__3389\ : IoSpan4Mux
    port map (
            O => \N__16435\,
            I => \N__16426\
        );

    \I__3388\ : Span4Mux_h
    port map (
            O => \N__16432\,
            I => \N__16423\
        );

    \I__3387\ : Span4Mux_v
    port map (
            O => \N__16429\,
            I => \N__16420\
        );

    \I__3386\ : Span4Mux_s3_h
    port map (
            O => \N__16426\,
            I => \N__16417\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__16423\,
            I => \resetGen_rst_1_iso\
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__16420\,
            I => \resetGen_rst_1_iso\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__16417\,
            I => \resetGen_rst_1_iso\
        );

    \I__3382\ : CEMux
    port map (
            O => \N__16410\,
            I => \N__16407\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__16407\,
            I => \N__16404\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__16404\,
            I => \N__16401\
        );

    \I__3379\ : Span4Mux_v
    port map (
            O => \N__16401\,
            I => \N__16398\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__16398\,
            I => \Lab_UT.scdp.u0.sccDnibble1En_0\
        );

    \I__3377\ : InMux
    port map (
            O => \N__16395\,
            I => \N__16392\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16392\,
            I => \N__16389\
        );

    \I__3375\ : Span4Mux_s3_h
    port map (
            O => \N__16389\,
            I => \N__16386\
        );

    \I__3374\ : Span4Mux_h
    port map (
            O => \N__16386\,
            I => \N__16383\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__16383\,
            I => \Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0dup_1\
        );

    \I__3372\ : InMux
    port map (
            O => \N__16380\,
            I => \N__16377\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__16377\,
            I => \Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__16374\,
            I => \Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93_cascade_\
        );

    \I__3369\ : SRMux
    port map (
            O => \N__16371\,
            I => \N__16368\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__16368\,
            I => \Lab_UT.scctrl.N_69_i\
        );

    \I__3367\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16362\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__16362\,
            I => \Lab_UT.scctrl.N_11\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__16359\,
            I => \N__16355\
        );

    \I__3364\ : InMux
    port map (
            O => \N__16358\,
            I => \N__16349\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16340\
        );

    \I__3362\ : InMux
    port map (
            O => \N__16354\,
            I => \N__16340\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16353\,
            I => \N__16340\
        );

    \I__3360\ : InMux
    port map (
            O => \N__16352\,
            I => \N__16340\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__16349\,
            I => \N__16337\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__16340\,
            I => \Lab_UT.scctrl.next_state_rst\
        );

    \I__3357\ : Odrv4
    port map (
            O => \N__16337\,
            I => \Lab_UT.scctrl.next_state_rst\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__16332\,
            I => \Lab_UT.scctrl.g0_9_a2_5_cascade_\
        );

    \I__3355\ : InMux
    port map (
            O => \N__16329\,
            I => \N__16323\
        );

    \I__3354\ : InMux
    port map (
            O => \N__16328\,
            I => \N__16323\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16323\,
            I => \Lab_UT.scctrl.next_state_rst_0_3_tz\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__16320\,
            I => \Lab_UT.scctrl.next_state_rst_0_3_0_cascade_\
        );

    \I__3351\ : InMux
    port map (
            O => \N__16317\,
            I => \N__16313\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__16316\,
            I => \N__16310\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__16313\,
            I => \N__16307\
        );

    \I__3348\ : InMux
    port map (
            O => \N__16310\,
            I => \N__16302\
        );

    \I__3347\ : Span4Mux_v
    port map (
            O => \N__16307\,
            I => \N__16299\
        );

    \I__3346\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16296\
        );

    \I__3345\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16293\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__16302\,
            I => \N__16288\
        );

    \I__3343\ : Span4Mux_s2_h
    port map (
            O => \N__16299\,
            I => \N__16288\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__16296\,
            I => rst_i_fast
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__16293\,
            I => rst_i_fast
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__16288\,
            I => rst_i_fast
        );

    \I__3339\ : InMux
    port map (
            O => \N__16281\,
            I => \N__16276\
        );

    \I__3338\ : InMux
    port map (
            O => \N__16280\,
            I => \N__16273\
        );

    \I__3337\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16270\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__16276\,
            I => \N__16267\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__16273\,
            I => \N__16264\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__16270\,
            I => \Lab_UT.scctrl.state_fast_3\
        );

    \I__3333\ : Odrv12
    port map (
            O => \N__16267\,
            I => \Lab_UT.scctrl.state_fast_3\
        );

    \I__3332\ : Odrv4
    port map (
            O => \N__16264\,
            I => \Lab_UT.scctrl.state_fast_3\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__16257\,
            I => \Lab_UT.scctrl.g0_0_0_0_cascade_\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__16254\,
            I => \Lab_UT.scctrl.g0_0_2_cascade_\
        );

    \I__3329\ : InMux
    port map (
            O => \N__16251\,
            I => \N__16248\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__16248\,
            I => \Lab_UT.scctrl.g0_0_3\
        );

    \I__3327\ : InMux
    port map (
            O => \N__16245\,
            I => \N__16242\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__16242\,
            I => \N__16238\
        );

    \I__3325\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16235\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__16238\,
            I => \buart__rx_shifter_1_fast_0\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__16235\,
            I => \buart__rx_shifter_1_fast_0\
        );

    \I__3322\ : InMux
    port map (
            O => \N__16230\,
            I => \N__16227\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__16227\,
            I => \Lab_UT.scctrl.N_408_0\
        );

    \I__3320\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16221\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__16221\,
            I => \Lab_UT.scctrl.g2_0_0\
        );

    \I__3318\ : InMux
    port map (
            O => \N__16218\,
            I => \N__16215\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__16215\,
            I => \Lab_UT.scctrl.N_17\
        );

    \I__3316\ : InMux
    port map (
            O => \N__16212\,
            I => \N__16201\
        );

    \I__3315\ : InMux
    port map (
            O => \N__16211\,
            I => \N__16201\
        );

    \I__3314\ : InMux
    port map (
            O => \N__16210\,
            I => \N__16198\
        );

    \I__3313\ : InMux
    port map (
            O => \N__16209\,
            I => \N__16193\
        );

    \I__3312\ : InMux
    port map (
            O => \N__16208\,
            I => \N__16193\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16207\,
            I => \N__16186\
        );

    \I__3310\ : InMux
    port map (
            O => \N__16206\,
            I => \N__16186\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__16201\,
            I => \N__16183\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__16198\,
            I => \N__16178\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__16193\,
            I => \N__16178\
        );

    \I__3306\ : InMux
    port map (
            O => \N__16192\,
            I => \N__16173\
        );

    \I__3305\ : InMux
    port map (
            O => \N__16191\,
            I => \N__16173\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__16186\,
            I => \Lab_UT.scctrl.N_240_i_0\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__16183\,
            I => \Lab_UT.scctrl.N_240_i_0\
        );

    \I__3302\ : Odrv12
    port map (
            O => \N__16178\,
            I => \Lab_UT.scctrl.N_240_i_0\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__16173\,
            I => \Lab_UT.scctrl.N_240_i_0\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__16164\,
            I => \N__16159\
        );

    \I__3299\ : InMux
    port map (
            O => \N__16163\,
            I => \N__16139\
        );

    \I__3298\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16139\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16139\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16158\,
            I => \N__16135\
        );

    \I__3295\ : InMux
    port map (
            O => \N__16157\,
            I => \N__16132\
        );

    \I__3294\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16121\
        );

    \I__3293\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16121\
        );

    \I__3292\ : InMux
    port map (
            O => \N__16154\,
            I => \N__16121\
        );

    \I__3291\ : InMux
    port map (
            O => \N__16153\,
            I => \N__16121\
        );

    \I__3290\ : InMux
    port map (
            O => \N__16152\,
            I => \N__16121\
        );

    \I__3289\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16118\
        );

    \I__3288\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16113\
        );

    \I__3287\ : InMux
    port map (
            O => \N__16149\,
            I => \N__16113\
        );

    \I__3286\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16108\
        );

    \I__3285\ : InMux
    port map (
            O => \N__16147\,
            I => \N__16108\
        );

    \I__3284\ : CascadeMux
    port map (
            O => \N__16146\,
            I => \N__16105\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__16139\,
            I => \N__16101\
        );

    \I__3282\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16096\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__16135\,
            I => \N__16093\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__16132\,
            I => \N__16088\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__16121\,
            I => \N__16088\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__16118\,
            I => \N__16081\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__16113\,
            I => \N__16081\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__16108\,
            I => \N__16081\
        );

    \I__3275\ : InMux
    port map (
            O => \N__16105\,
            I => \N__16078\
        );

    \I__3274\ : InMux
    port map (
            O => \N__16104\,
            I => \N__16075\
        );

    \I__3273\ : Span4Mux_v
    port map (
            O => \N__16101\,
            I => \N__16072\
        );

    \I__3272\ : InMux
    port map (
            O => \N__16100\,
            I => \N__16067\
        );

    \I__3271\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16067\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__16096\,
            I => \N__16056\
        );

    \I__3269\ : Span4Mux_v
    port map (
            O => \N__16093\,
            I => \N__16056\
        );

    \I__3268\ : Span4Mux_v
    port map (
            O => \N__16088\,
            I => \N__16056\
        );

    \I__3267\ : Span4Mux_v
    port map (
            O => \N__16081\,
            I => \N__16056\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__16078\,
            I => \N__16056\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__16075\,
            I => \N__16051\
        );

    \I__3264\ : Span4Mux_s2_h
    port map (
            O => \N__16072\,
            I => \N__16051\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__16067\,
            I => bu_rx_data_i_1_5
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__16056\,
            I => bu_rx_data_i_1_5
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__16051\,
            I => bu_rx_data_i_1_5
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__16044\,
            I => \Lab_UT.scctrl.N_412_cascade_\
        );

    \I__3259\ : InMux
    port map (
            O => \N__16041\,
            I => \N__16035\
        );

    \I__3258\ : InMux
    port map (
            O => \N__16040\,
            I => \N__16035\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__16035\,
            I => \Lab_UT.scctrl.next_state_rst_0_1\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__16032\,
            I => \Lab_UT.scctrl.state_ret_4_RNOZ0Z_10_cascade_\
        );

    \I__3255\ : InMux
    port map (
            O => \N__16029\,
            I => \N__16026\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__16026\,
            I => \N__16023\
        );

    \I__3253\ : Span4Mux_v
    port map (
            O => \N__16023\,
            I => \N__16020\
        );

    \I__3252\ : Odrv4
    port map (
            O => \N__16020\,
            I => \Lab_UT.scctrl.state_ret_4_RNOZ0Z_6\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__16017\,
            I => \N__16014\
        );

    \I__3250\ : InMux
    port map (
            O => \N__16014\,
            I => \N__16007\
        );

    \I__3249\ : InMux
    port map (
            O => \N__16013\,
            I => \N__16007\
        );

    \I__3248\ : InMux
    port map (
            O => \N__16012\,
            I => \N__16004\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__16007\,
            I => \N__15999\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__16004\,
            I => \N__15999\
        );

    \I__3245\ : Span4Mux_v
    port map (
            O => \N__15999\,
            I => \N__15996\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__15996\,
            I => \Lab_UT.scctrl.N_295\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__15993\,
            I => \Lab_UT.scctrl.N_295_cascade_\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15987\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__15987\,
            I => \N__15984\
        );

    \I__3240\ : Sp12to4
    port map (
            O => \N__15984\,
            I => \N__15981\
        );

    \I__3239\ : Odrv12
    port map (
            O => \N__15981\,
            I => \Lab_UT.scctrl.N_40_i\
        );

    \I__3238\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15971\
        );

    \I__3237\ : CascadeMux
    port map (
            O => \N__15977\,
            I => \N__15968\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__15976\,
            I => \N__15965\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__15975\,
            I => \N__15962\
        );

    \I__3234\ : CascadeMux
    port map (
            O => \N__15974\,
            I => \N__15959\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__15971\,
            I => \N__15956\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15968\,
            I => \N__15953\
        );

    \I__3231\ : InMux
    port map (
            O => \N__15965\,
            I => \N__15949\
        );

    \I__3230\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15944\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15944\
        );

    \I__3228\ : Span4Mux_h
    port map (
            O => \N__15956\,
            I => \N__15941\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__15953\,
            I => \N__15938\
        );

    \I__3226\ : InMux
    port map (
            O => \N__15952\,
            I => \N__15935\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__15949\,
            I => \Lab_UT.scctrl.N_487\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15944\,
            I => \Lab_UT.scctrl.N_487\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__15941\,
            I => \Lab_UT.scctrl.N_487\
        );

    \I__3222\ : Odrv4
    port map (
            O => \N__15938\,
            I => \Lab_UT.scctrl.N_487\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__15935\,
            I => \Lab_UT.scctrl.N_487\
        );

    \I__3220\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15921\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__15921\,
            I => \N__15916\
        );

    \I__3218\ : InMux
    port map (
            O => \N__15920\,
            I => \N__15911\
        );

    \I__3217\ : InMux
    port map (
            O => \N__15919\,
            I => \N__15911\
        );

    \I__3216\ : Span4Mux_h
    port map (
            O => \N__15916\,
            I => \N__15908\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__15911\,
            I => \Lab_UT.scctrl.N_284\
        );

    \I__3214\ : Odrv4
    port map (
            O => \N__15908\,
            I => \Lab_UT.scctrl.N_284\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__15903\,
            I => \N__15897\
        );

    \I__3212\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15893\
        );

    \I__3211\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15888\
        );

    \I__3210\ : InMux
    port map (
            O => \N__15900\,
            I => \N__15885\
        );

    \I__3209\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15880\
        );

    \I__3208\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15880\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__15893\,
            I => \N__15875\
        );

    \I__3206\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15870\
        );

    \I__3205\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15870\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__15888\,
            I => \N__15865\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__15885\,
            I => \N__15865\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__15880\,
            I => \N__15862\
        );

    \I__3201\ : InMux
    port map (
            O => \N__15879\,
            I => \N__15859\
        );

    \I__3200\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15856\
        );

    \I__3199\ : Span4Mux_v
    port map (
            O => \N__15875\,
            I => \N__15853\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__15870\,
            I => \N__15842\
        );

    \I__3197\ : Span4Mux_v
    port map (
            O => \N__15865\,
            I => \N__15842\
        );

    \I__3196\ : Span4Mux_v
    port map (
            O => \N__15862\,
            I => \N__15842\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__15859\,
            I => \N__15842\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__15856\,
            I => \N__15842\
        );

    \I__3193\ : Odrv4
    port map (
            O => \N__15853\,
            I => \Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__15842\,
            I => \Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__15837\,
            I => \Lab_UT.scctrl.N_408_cascade_\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__15834\,
            I => \Lab_UT.scctrl.g0_i_a8_0_1_cascade_\
        );

    \I__3189\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15828\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__15828\,
            I => \N__15825\
        );

    \I__3187\ : Span4Mux_h
    port map (
            O => \N__15825\,
            I => \N__15822\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__15822\,
            I => \Lab_UT.scctrl.G_24_i_o7_0_0\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__15819\,
            I => \Lab_UT.scctrl.N_12_1_cascade_\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__15816\,
            I => \N__15813\
        );

    \I__3183\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15810\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__15810\,
            I => \Lab_UT.scctrl.N_408\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__15807\,
            I => \Lab_UT.scctrl.N_418_2_cascade_\
        );

    \I__3180\ : InMux
    port map (
            O => \N__15804\,
            I => \N__15801\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__15801\,
            I => \N__15798\
        );

    \I__3178\ : Span4Mux_h
    port map (
            O => \N__15798\,
            I => \N__15795\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__15795\,
            I => \Lab_UT.scctrl.g1_0\
        );

    \I__3176\ : InMux
    port map (
            O => \N__15792\,
            I => \N__15784\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15791\,
            I => \N__15773\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15773\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15773\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15773\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15787\,
            I => \N__15773\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__15784\,
            I => \N__15770\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__15773\,
            I => \Lab_UT.scctrl.N_418\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__15770\,
            I => \Lab_UT.scctrl.N_418\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__15765\,
            I => \N__15761\
        );

    \I__3166\ : InMux
    port map (
            O => \N__15764\,
            I => \N__15756\
        );

    \I__3165\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15756\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__15756\,
            I => \N__15753\
        );

    \I__3163\ : Span4Mux_s3_h
    port map (
            O => \N__15753\,
            I => \N__15750\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__15750\,
            I => \Lab_UT.scctrl.N_415\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15747\,
            I => \N__15744\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__15744\,
            I => \N__15738\
        );

    \I__3159\ : InMux
    port map (
            O => \N__15743\,
            I => \N__15735\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15742\,
            I => \N__15730\
        );

    \I__3157\ : InMux
    port map (
            O => \N__15741\,
            I => \N__15730\
        );

    \I__3156\ : Span4Mux_s2_v
    port map (
            O => \N__15738\,
            I => \N__15727\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__15735\,
            I => \Lab_UT.scctrl.state_ret_0_fastZ0\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__15730\,
            I => \Lab_UT.scctrl.state_ret_0_fastZ0\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__15727\,
            I => \Lab_UT.scctrl.state_ret_0_fastZ0\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__15720\,
            I => \Lab_UT.scctrl.next_state_rst_4_4_cascade_\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15717\,
            I => \N__15714\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__15714\,
            I => \Lab_UT.scctrl.N_290_1\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__15711\,
            I => \N__15708\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15708\,
            I => \N__15705\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__15705\,
            I => \Lab_UT.scctrl.g0_1_0\
        );

    \I__3146\ : InMux
    port map (
            O => \N__15702\,
            I => \N__15699\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__15699\,
            I => \N__15692\
        );

    \I__3144\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15685\
        );

    \I__3143\ : InMux
    port map (
            O => \N__15697\,
            I => \N__15685\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15696\,
            I => \N__15685\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15695\,
            I => \N__15682\
        );

    \I__3140\ : Span4Mux_v
    port map (
            O => \N__15692\,
            I => \N__15679\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__15685\,
            I => \Lab_UT.scctrl.next_state_rst_1_3\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__15682\,
            I => \Lab_UT.scctrl.next_state_rst_1_3\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__15679\,
            I => \Lab_UT.scctrl.next_state_rst_1_3\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__15672\,
            I => \Lab_UT.scctrl.next_state_rst_4_2_cascade_\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15669\,
            I => \N__15666\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__15666\,
            I => \Lab_UT.scctrl.N_290\
        );

    \I__3133\ : InMux
    port map (
            O => \N__15663\,
            I => \N__15660\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__15660\,
            I => \N__15657\
        );

    \I__3131\ : Odrv4
    port map (
            O => \N__15657\,
            I => \Lab_UT.scctrl.next_state_0_3\
        );

    \I__3130\ : InMux
    port map (
            O => \N__15654\,
            I => \N__15651\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__15651\,
            I => \Lab_UT.scctrl.N_415_2\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__15648\,
            I => \Lab_UT.scctrl.g1_2_0_cascade_\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__15645\,
            I => \Lab_UT.scctrl.next_stateZ0Z_2_cascade_\
        );

    \I__3126\ : InMux
    port map (
            O => \N__15642\,
            I => \N__15636\
        );

    \I__3125\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15636\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__15636\,
            I => \N__15633\
        );

    \I__3123\ : Span4Mux_h
    port map (
            O => \N__15633\,
            I => \N__15630\
        );

    \I__3122\ : Span4Mux_v
    port map (
            O => \N__15630\,
            I => \N__15627\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__15627\,
            I => \Lab_UT.scctrl.next_state_rst_2\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__15624\,
            I => \N__15621\
        );

    \I__3119\ : InMux
    port map (
            O => \N__15621\,
            I => \N__15617\
        );

    \I__3118\ : InMux
    port map (
            O => \N__15620\,
            I => \N__15614\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__15617\,
            I => \N__15608\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__15614\,
            I => \N__15608\
        );

    \I__3115\ : InMux
    port map (
            O => \N__15613\,
            I => \N__15605\
        );

    \I__3114\ : Span4Mux_v
    port map (
            O => \N__15608\,
            I => \N__15602\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__15605\,
            I => \Lab_UT.scctrl.next_stateZ0Z_2\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__15602\,
            I => \Lab_UT.scctrl.next_stateZ0Z_2\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__15597\,
            I => \N__15593\
        );

    \I__3110\ : CascadeMux
    port map (
            O => \N__15596\,
            I => \N__15590\
        );

    \I__3109\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15576\
        );

    \I__3108\ : InMux
    port map (
            O => \N__15590\,
            I => \N__15576\
        );

    \I__3107\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15576\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15588\,
            I => \N__15576\
        );

    \I__3105\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15576\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__15576\,
            I => \N__15573\
        );

    \I__3103\ : Odrv4
    port map (
            O => \N__15573\,
            I => \Lab_UT.scctrl.g1_1_1_0\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15570\,
            I => \N__15558\
        );

    \I__3101\ : InMux
    port map (
            O => \N__15569\,
            I => \N__15558\
        );

    \I__3100\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15558\
        );

    \I__3099\ : InMux
    port map (
            O => \N__15567\,
            I => \N__15558\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__15558\,
            I => \Lab_UT.scctrl.g1_2_0\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__15555\,
            I => \Lab_UT.scctrl.next_state_rst_4_3_cascade_\
        );

    \I__3096\ : InMux
    port map (
            O => \N__15552\,
            I => \N__15549\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15549\,
            I => \N__15546\
        );

    \I__3094\ : Odrv4
    port map (
            O => \N__15546\,
            I => \Lab_UT.scctrl.N_290_0\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15543\,
            I => \N__15540\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__15540\,
            I => \Lab_UT.scctrl.next_state_rst_4_5\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__15537\,
            I => \Lab_UT.scctrl.N_20_i_cascade_\
        );

    \I__3090\ : InMux
    port map (
            O => \N__15534\,
            I => \N__15531\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__15531\,
            I => \Lab_UT.scctrl.N_277\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__15528\,
            I => \Lab_UT.scctrl.N_277_cascade_\
        );

    \I__3087\ : IoInMux
    port map (
            O => \N__15525\,
            I => \N__15522\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__15522\,
            I => \N__15519\
        );

    \I__3085\ : IoSpan4Mux
    port map (
            O => \N__15519\,
            I => \N__15516\
        );

    \I__3084\ : Span4Mux_s3_h
    port map (
            O => \N__15516\,
            I => \N__15513\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__15513\,
            I => \N_67\
        );

    \I__3082\ : InMux
    port map (
            O => \N__15510\,
            I => \N__15507\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__15507\,
            I => \Lab_UT.scctrl.N_355\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15504\,
            I => \N__15500\
        );

    \I__3079\ : InMux
    port map (
            O => \N__15503\,
            I => \N__15491\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__15500\,
            I => \N__15488\
        );

    \I__3077\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15479\
        );

    \I__3076\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15479\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15479\
        );

    \I__3074\ : InMux
    port map (
            O => \N__15496\,
            I => \N__15479\
        );

    \I__3073\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15474\
        );

    \I__3072\ : InMux
    port map (
            O => \N__15494\,
            I => \N__15474\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__15491\,
            I => \Lab_UT.scctrl.N_36\
        );

    \I__3070\ : Odrv4
    port map (
            O => \N__15488\,
            I => \Lab_UT.scctrl.N_36\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__15479\,
            I => \Lab_UT.scctrl.N_36\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__15474\,
            I => \Lab_UT.scctrl.N_36\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__15465\,
            I => \Lab_UT.scctrl.N_27_i_cascade_\
        );

    \I__3066\ : InMux
    port map (
            O => \N__15462\,
            I => \N__15452\
        );

    \I__3065\ : InMux
    port map (
            O => \N__15461\,
            I => \N__15444\
        );

    \I__3064\ : InMux
    port map (
            O => \N__15460\,
            I => \N__15440\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15459\,
            I => \N__15437\
        );

    \I__3062\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15434\
        );

    \I__3061\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15431\
        );

    \I__3060\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15425\
        );

    \I__3059\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15425\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__15452\,
            I => \N__15422\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15419\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15450\,
            I => \N__15416\
        );

    \I__3055\ : InMux
    port map (
            O => \N__15449\,
            I => \N__15411\
        );

    \I__3054\ : InMux
    port map (
            O => \N__15448\,
            I => \N__15411\
        );

    \I__3053\ : InMux
    port map (
            O => \N__15447\,
            I => \N__15408\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__15444\,
            I => \N__15405\
        );

    \I__3051\ : InMux
    port map (
            O => \N__15443\,
            I => \N__15402\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__15440\,
            I => \N__15399\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__15437\,
            I => \N__15395\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__15434\,
            I => \N__15390\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__15431\,
            I => \N__15390\
        );

    \I__3046\ : CascadeMux
    port map (
            O => \N__15430\,
            I => \N__15387\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__15425\,
            I => \N__15380\
        );

    \I__3044\ : Span4Mux_h
    port map (
            O => \N__15422\,
            I => \N__15380\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__15419\,
            I => \N__15380\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__15416\,
            I => \N__15377\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__15411\,
            I => \N__15374\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15408\,
            I => \N__15367\
        );

    \I__3039\ : Span4Mux_v
    port map (
            O => \N__15405\,
            I => \N__15367\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__15402\,
            I => \N__15367\
        );

    \I__3037\ : Span4Mux_h
    port map (
            O => \N__15399\,
            I => \N__15364\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15361\
        );

    \I__3035\ : Span4Mux_v
    port map (
            O => \N__15395\,
            I => \N__15358\
        );

    \I__3034\ : Span4Mux_h
    port map (
            O => \N__15390\,
            I => \N__15355\
        );

    \I__3033\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15352\
        );

    \I__3032\ : Span4Mux_v
    port map (
            O => \N__15380\,
            I => \N__15347\
        );

    \I__3031\ : Span4Mux_v
    port map (
            O => \N__15377\,
            I => \N__15347\
        );

    \I__3030\ : Span4Mux_s3_h
    port map (
            O => \N__15374\,
            I => \N__15340\
        );

    \I__3029\ : Span4Mux_h
    port map (
            O => \N__15367\,
            I => \N__15340\
        );

    \I__3028\ : Span4Mux_v
    port map (
            O => \N__15364\,
            I => \N__15340\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__15361\,
            I => rst_i
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__15358\,
            I => rst_i
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__15355\,
            I => rst_i
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__15352\,
            I => rst_i
        );

    \I__3023\ : Odrv4
    port map (
            O => \N__15347\,
            I => rst_i
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__15340\,
            I => rst_i
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__15327\,
            I => \N__15324\
        );

    \I__3020\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15321\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__15321\,
            I => \Lab_UT.scctrl.N_19\
        );

    \I__3018\ : InMux
    port map (
            O => \N__15318\,
            I => \N__15315\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__15315\,
            I => \Lab_UT.scctrl.G_24_i_1_0\
        );

    \I__3016\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15308\
        );

    \I__3015\ : InMux
    port map (
            O => \N__15311\,
            I => \N__15305\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__15308\,
            I => \N__15302\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__15305\,
            I => \N__15299\
        );

    \I__3012\ : Span4Mux_h
    port map (
            O => \N__15302\,
            I => \N__15296\
        );

    \I__3011\ : Odrv12
    port map (
            O => \N__15299\,
            I => \Lab_UT.scctrl.N_401_0\
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__15296\,
            I => \Lab_UT.scctrl.N_401_0\
        );

    \I__3009\ : InMux
    port map (
            O => \N__15291\,
            I => \N__15288\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__15288\,
            I => \N__15284\
        );

    \I__3007\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15281\
        );

    \I__3006\ : Span4Mux_h
    port map (
            O => \N__15284\,
            I => \N__15278\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__15281\,
            I => \N__15275\
        );

    \I__3004\ : Span4Mux_v
    port map (
            O => \N__15278\,
            I => \N__15272\
        );

    \I__3003\ : Span4Mux_h
    port map (
            O => \N__15275\,
            I => \N__15269\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__15272\,
            I => \Lab_UT.scctrl.N_9_0\
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__15269\,
            I => \Lab_UT.scctrl.N_9_0\
        );

    \I__3000\ : InMux
    port map (
            O => \N__15264\,
            I => \N__15261\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__15261\,
            I => \N__15258\
        );

    \I__2998\ : Span4Mux_v
    port map (
            O => \N__15258\,
            I => \N__15254\
        );

    \I__2997\ : InMux
    port map (
            O => \N__15257\,
            I => \N__15251\
        );

    \I__2996\ : Odrv4
    port map (
            O => \N__15254\,
            I => \Lab_UT.scctrl.g0_i_2\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__15251\,
            I => \Lab_UT.scctrl.g0_i_2\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__15246\,
            I => \Lab_UT.scctrl.N_170_i_cascade_\
        );

    \I__2993\ : InMux
    port map (
            O => \N__15243\,
            I => \N__15240\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__15240\,
            I => \Lab_UT.scctrl.G_24_i_o6_0_0\
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__15237\,
            I => \Lab_UT.scctrl.N_17_i_cascade_\
        );

    \I__2990\ : InMux
    port map (
            O => \N__15234\,
            I => \N__15231\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__15231\,
            I => \Lab_UT.scctrl.N_418_1\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__15228\,
            I => \Lab_UT.scctrl.g0_8_0_cascade_\
        );

    \I__2987\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15222\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__15222\,
            I => \Lab_UT.scctrl.g0_8_2\
        );

    \I__2985\ : CascadeMux
    port map (
            O => \N__15219\,
            I => \N__15215\
        );

    \I__2984\ : InMux
    port map (
            O => \N__15218\,
            I => \N__15210\
        );

    \I__2983\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15210\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__15210\,
            I => \N__15207\
        );

    \I__2981\ : Span4Mux_v
    port map (
            O => \N__15207\,
            I => \N__15204\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__15204\,
            I => \Lab_UT.scctrl.N_444_1\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__15201\,
            I => \N__15198\
        );

    \I__2978\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15190\
        );

    \I__2977\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15190\
        );

    \I__2976\ : InMux
    port map (
            O => \N__15196\,
            I => \N__15187\
        );

    \I__2975\ : InMux
    port map (
            O => \N__15195\,
            I => \N__15184\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__15190\,
            I => \N__15177\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__15187\,
            I => \N__15172\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__15184\,
            I => \N__15172\
        );

    \I__2971\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15165\
        );

    \I__2970\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15162\
        );

    \I__2969\ : InMux
    port map (
            O => \N__15181\,
            I => \N__15159\
        );

    \I__2968\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15156\
        );

    \I__2967\ : Span4Mux_v
    port map (
            O => \N__15177\,
            I => \N__15151\
        );

    \I__2966\ : Span4Mux_v
    port map (
            O => \N__15172\,
            I => \N__15151\
        );

    \I__2965\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15142\
        );

    \I__2964\ : InMux
    port map (
            O => \N__15170\,
            I => \N__15142\
        );

    \I__2963\ : InMux
    port map (
            O => \N__15169\,
            I => \N__15142\
        );

    \I__2962\ : InMux
    port map (
            O => \N__15168\,
            I => \N__15142\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__15165\,
            I => bu_rx_data_i_1_6
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__15162\,
            I => bu_rx_data_i_1_6
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__15159\,
            I => bu_rx_data_i_1_6
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__15156\,
            I => bu_rx_data_i_1_6
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__15151\,
            I => bu_rx_data_i_1_6
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__15142\,
            I => bu_rx_data_i_1_6
        );

    \I__2955\ : InMux
    port map (
            O => \N__15129\,
            I => \N__15121\
        );

    \I__2954\ : InMux
    port map (
            O => \N__15128\,
            I => \N__15117\
        );

    \I__2953\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15113\
        );

    \I__2952\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15108\
        );

    \I__2951\ : InMux
    port map (
            O => \N__15125\,
            I => \N__15108\
        );

    \I__2950\ : InMux
    port map (
            O => \N__15124\,
            I => \N__15101\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__15121\,
            I => \N__15098\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__15120\,
            I => \N__15093\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__15117\,
            I => \N__15088\
        );

    \I__2946\ : InMux
    port map (
            O => \N__15116\,
            I => \N__15085\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__15113\,
            I => \N__15080\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__15108\,
            I => \N__15076\
        );

    \I__2943\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15064\
        );

    \I__2942\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15064\
        );

    \I__2941\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15061\
        );

    \I__2940\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15058\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__15101\,
            I => \N__15053\
        );

    \I__2938\ : Span4Mux_h
    port map (
            O => \N__15098\,
            I => \N__15053\
        );

    \I__2937\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15042\
        );

    \I__2936\ : InMux
    port map (
            O => \N__15096\,
            I => \N__15042\
        );

    \I__2935\ : InMux
    port map (
            O => \N__15093\,
            I => \N__15042\
        );

    \I__2934\ : InMux
    port map (
            O => \N__15092\,
            I => \N__15042\
        );

    \I__2933\ : InMux
    port map (
            O => \N__15091\,
            I => \N__15042\
        );

    \I__2932\ : Span12Mux_s5_h
    port map (
            O => \N__15088\,
            I => \N__15039\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__15085\,
            I => \N__15036\
        );

    \I__2930\ : InMux
    port map (
            O => \N__15084\,
            I => \N__15033\
        );

    \I__2929\ : InMux
    port map (
            O => \N__15083\,
            I => \N__15030\
        );

    \I__2928\ : Span4Mux_v
    port map (
            O => \N__15080\,
            I => \N__15027\
        );

    \I__2927\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15024\
        );

    \I__2926\ : Span4Mux_v
    port map (
            O => \N__15076\,
            I => \N__15021\
        );

    \I__2925\ : InMux
    port map (
            O => \N__15075\,
            I => \N__15018\
        );

    \I__2924\ : InMux
    port map (
            O => \N__15074\,
            I => \N__15009\
        );

    \I__2923\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15009\
        );

    \I__2922\ : InMux
    port map (
            O => \N__15072\,
            I => \N__15009\
        );

    \I__2921\ : InMux
    port map (
            O => \N__15071\,
            I => \N__15009\
        );

    \I__2920\ : InMux
    port map (
            O => \N__15070\,
            I => \N__15004\
        );

    \I__2919\ : InMux
    port map (
            O => \N__15069\,
            I => \N__15004\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__15064\,
            I => \N__14999\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__15061\,
            I => \N__14999\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__15058\,
            I => \N__14994\
        );

    \I__2915\ : Span4Mux_v
    port map (
            O => \N__15053\,
            I => \N__14994\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__15042\,
            I => \N__14991\
        );

    \I__2913\ : Odrv12
    port map (
            O => \N__15039\,
            I => bu_rx_data_4
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__15036\,
            I => bu_rx_data_4
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__15033\,
            I => bu_rx_data_4
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__15030\,
            I => bu_rx_data_4
        );

    \I__2909\ : Odrv4
    port map (
            O => \N__15027\,
            I => bu_rx_data_4
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__15024\,
            I => bu_rx_data_4
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__15021\,
            I => bu_rx_data_4
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__15018\,
            I => bu_rx_data_4
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__15009\,
            I => bu_rx_data_4
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__15004\,
            I => bu_rx_data_4
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__14999\,
            I => bu_rx_data_4
        );

    \I__2902\ : Odrv4
    port map (
            O => \N__14994\,
            I => bu_rx_data_4
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__14991\,
            I => bu_rx_data_4
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__14964\,
            I => \Lab_UT.scctrl.G_24_i_a6_2_2_cascade_\
        );

    \I__2899\ : InMux
    port map (
            O => \N__14961\,
            I => \N__14958\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__14958\,
            I => \N__14955\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__14955\,
            I => \N__14952\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__14952\,
            I => \Lab_UT.scctrl.N_12_3\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__14949\,
            I => \N__14945\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__14948\,
            I => \N__14942\
        );

    \I__2893\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14932\
        );

    \I__2892\ : InMux
    port map (
            O => \N__14942\,
            I => \N__14927\
        );

    \I__2891\ : InMux
    port map (
            O => \N__14941\,
            I => \N__14927\
        );

    \I__2890\ : InMux
    port map (
            O => \N__14940\,
            I => \N__14923\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__14939\,
            I => \N__14920\
        );

    \I__2888\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14913\
        );

    \I__2887\ : InMux
    port map (
            O => \N__14937\,
            I => \N__14913\
        );

    \I__2886\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14913\
        );

    \I__2885\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14910\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__14932\,
            I => \N__14904\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__14927\,
            I => \N__14904\
        );

    \I__2882\ : InMux
    port map (
            O => \N__14926\,
            I => \N__14901\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__14923\,
            I => \N__14897\
        );

    \I__2880\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14894\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__14913\,
            I => \N__14891\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__14910\,
            I => \N__14888\
        );

    \I__2877\ : InMux
    port map (
            O => \N__14909\,
            I => \N__14885\
        );

    \I__2876\ : Span4Mux_h
    port map (
            O => \N__14904\,
            I => \N__14882\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__14901\,
            I => \N__14879\
        );

    \I__2874\ : InMux
    port map (
            O => \N__14900\,
            I => \N__14876\
        );

    \I__2873\ : Span12Mux_s11_v
    port map (
            O => \N__14897\,
            I => \N__14871\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__14894\,
            I => \N__14871\
        );

    \I__2871\ : Span4Mux_h
    port map (
            O => \N__14891\,
            I => \N__14860\
        );

    \I__2870\ : Span4Mux_h
    port map (
            O => \N__14888\,
            I => \N__14860\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__14885\,
            I => \N__14860\
        );

    \I__2868\ : Span4Mux_v
    port map (
            O => \N__14882\,
            I => \N__14860\
        );

    \I__2867\ : Span4Mux_h
    port map (
            O => \N__14879\,
            I => \N__14860\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__14876\,
            I => bu_rx_data_6
        );

    \I__2865\ : Odrv12
    port map (
            O => \N__14871\,
            I => bu_rx_data_6
        );

    \I__2864\ : Odrv4
    port map (
            O => \N__14860\,
            I => bu_rx_data_6
        );

    \I__2863\ : InMux
    port map (
            O => \N__14853\,
            I => \N__14843\
        );

    \I__2862\ : InMux
    port map (
            O => \N__14852\,
            I => \N__14843\
        );

    \I__2861\ : InMux
    port map (
            O => \N__14851\,
            I => \N__14843\
        );

    \I__2860\ : InMux
    port map (
            O => \N__14850\,
            I => \N__14840\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__14843\,
            I => \N__14837\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__14840\,
            I => \N__14833\
        );

    \I__2857\ : Span12Mux_s9_v
    port map (
            O => \N__14837\,
            I => \N__14830\
        );

    \I__2856\ : InMux
    port map (
            O => \N__14836\,
            I => \N__14827\
        );

    \I__2855\ : Odrv4
    port map (
            O => \N__14833\,
            I => \Lab_UT.scctrl.N_241_i_0\
        );

    \I__2854\ : Odrv12
    port map (
            O => \N__14830\,
            I => \Lab_UT.scctrl.N_241_i_0\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__14827\,
            I => \Lab_UT.scctrl.N_241_i_0\
        );

    \I__2852\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14817\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__14817\,
            I => \Lab_UT.scctrl.G_24_i_2_0\
        );

    \I__2850\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14811\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__14811\,
            I => \Lab_UT.scctrl.G_24_i_a6_0_2\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__14808\,
            I => \Lab_UT.scctrl.N_5_2_cascade_\
        );

    \I__2847\ : InMux
    port map (
            O => \N__14805\,
            I => \N__14802\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__14802\,
            I => \N__14799\
        );

    \I__2845\ : Odrv12
    port map (
            O => \N__14799\,
            I => \Lab_UT.scctrl.next_state_rst_2_1\
        );

    \I__2844\ : InMux
    port map (
            O => \N__14796\,
            I => \N__14793\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__14793\,
            I => \Lab_UT.scctrl.next_state_rst_4_1\
        );

    \I__2842\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14786\
        );

    \I__2841\ : InMux
    port map (
            O => \N__14789\,
            I => \N__14783\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__14786\,
            I => \Lab_UT.scctrl.G_15_0_a10_1_2\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__14783\,
            I => \Lab_UT.scctrl.G_15_0_a10_1_2\
        );

    \I__2838\ : InMux
    port map (
            O => \N__14778\,
            I => \N__14775\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__14775\,
            I => \Lab_UT.scctrl.N_7\
        );

    \I__2836\ : InMux
    port map (
            O => \N__14772\,
            I => \N__14769\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__14769\,
            I => \Lab_UT.scctrl.g0_8_0_0\
        );

    \I__2834\ : InMux
    port map (
            O => \N__14766\,
            I => \N__14763\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__14763\,
            I => \N__14759\
        );

    \I__2832\ : InMux
    port map (
            O => \N__14762\,
            I => \N__14756\
        );

    \I__2831\ : Span4Mux_v
    port map (
            O => \N__14759\,
            I => \N__14753\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__14756\,
            I => \N__14750\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__14753\,
            I => \Lab_UT.scctrl.N_223_0_0\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__14750\,
            I => \Lab_UT.scctrl.N_223_0_0\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__14745\,
            I => \Lab_UT.scctrl.N_419_0_cascade_\
        );

    \I__2826\ : InMux
    port map (
            O => \N__14742\,
            I => \N__14739\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14739\,
            I => \N__14736\
        );

    \I__2824\ : Span4Mux_h
    port map (
            O => \N__14736\,
            I => \N__14733\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__14733\,
            I => \Lab_UT.scctrl.g1\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__14730\,
            I => \N__14727\
        );

    \I__2821\ : InMux
    port map (
            O => \N__14727\,
            I => \N__14724\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__14724\,
            I => \N__14721\
        );

    \I__2819\ : Span4Mux_v
    port map (
            O => \N__14721\,
            I => \N__14718\
        );

    \I__2818\ : Odrv4
    port map (
            O => \N__14718\,
            I => \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_0_3\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__14715\,
            I => \Lab_UT.scctrl.g0_2_0_0_a3_2_cascade_\
        );

    \I__2816\ : InMux
    port map (
            O => \N__14712\,
            I => \N__14709\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__14709\,
            I => \N__14706\
        );

    \I__2814\ : Odrv12
    port map (
            O => \N__14706\,
            I => \Lab_UT.scctrl.G_24_i_a3_3\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__14703\,
            I => \Lab_UT.scctrl.G_24_i_a3_5_cascade_\
        );

    \I__2812\ : InMux
    port map (
            O => \N__14700\,
            I => \N__14697\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__14697\,
            I => \Lab_UT.scctrl.G_24_i_a3_0_3\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__14694\,
            I => \N__14691\
        );

    \I__2809\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14688\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__14688\,
            I => \Lab_UT.scctrl.G_24_i_a3_0_1\
        );

    \I__2807\ : InMux
    port map (
            O => \N__14685\,
            I => \N__14682\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__14682\,
            I => \N__14679\
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__14679\,
            I => \Lab_UT.scctrl.N_15\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__14676\,
            I => \N__14673\
        );

    \I__2803\ : InMux
    port map (
            O => \N__14673\,
            I => \N__14670\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__14670\,
            I => \Lab_UT.scctrl.next_state_rst_0_3_tz_0\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__14667\,
            I => \Lab_UT.scctrl.g0_0_4_cascade_\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__14664\,
            I => \Lab_UT.scctrl.next_state_rst_cascade_\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__14661\,
            I => \N__14657\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__14660\,
            I => \N__14654\
        );

    \I__2797\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14647\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14647\
        );

    \I__2795\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14644\
        );

    \I__2794\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14641\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__14647\,
            I => \N__14638\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__14644\,
            I => \N__14623\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14641\,
            I => \N__14623\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__14638\,
            I => \N__14623\
        );

    \I__2789\ : InMux
    port map (
            O => \N__14637\,
            I => \N__14612\
        );

    \I__2788\ : InMux
    port map (
            O => \N__14636\,
            I => \N__14612\
        );

    \I__2787\ : InMux
    port map (
            O => \N__14635\,
            I => \N__14612\
        );

    \I__2786\ : InMux
    port map (
            O => \N__14634\,
            I => \N__14612\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14633\,
            I => \N__14612\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14632\,
            I => \N__14609\
        );

    \I__2783\ : InMux
    port map (
            O => \N__14631\,
            I => \N__14604\
        );

    \I__2782\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14604\
        );

    \I__2781\ : Span4Mux_v
    port map (
            O => \N__14623\,
            I => \N__14599\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__14612\,
            I => \N__14599\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__14609\,
            I => \N__14596\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__14604\,
            I => \N__14593\
        );

    \I__2777\ : Span4Mux_v
    port map (
            O => \N__14599\,
            I => \N__14589\
        );

    \I__2776\ : Span4Mux_h
    port map (
            O => \N__14596\,
            I => \N__14584\
        );

    \I__2775\ : Span4Mux_v
    port map (
            O => \N__14593\,
            I => \N__14584\
        );

    \I__2774\ : InMux
    port map (
            O => \N__14592\,
            I => \N__14581\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__14589\,
            I => \Lab_UT.scctrl.state_i_1_0_rep2\
        );

    \I__2772\ : Odrv4
    port map (
            O => \N__14584\,
            I => \Lab_UT.scctrl.state_i_1_0_rep2\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__14581\,
            I => \Lab_UT.scctrl.state_i_1_0_rep2\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__14574\,
            I => \Lab_UT.scctrl.N_299_i_0_cascade_\
        );

    \I__2769\ : InMux
    port map (
            O => \N__14571\,
            I => \N__14567\
        );

    \I__2768\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14564\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__14567\,
            I => \N__14559\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__14564\,
            I => \N__14559\
        );

    \I__2765\ : Odrv4
    port map (
            O => \N__14559\,
            I => \Lab_UT.scctrl.N_4\
        );

    \I__2764\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14553\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__14553\,
            I => \Lab_UT.scctrl.N_240_reti\
        );

    \I__2762\ : InMux
    port map (
            O => \N__14550\,
            I => \N__14547\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__14547\,
            I => \Lab_UT.scctrl.N_419_1\
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__14544\,
            I => \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_2_3_cascade_\
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__14541\,
            I => \N__14538\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14538\,
            I => \N__14535\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__14535\,
            I => \N__14532\
        );

    \I__2756\ : Odrv4
    port map (
            O => \N__14532\,
            I => \Lab_UT.scctrl.g0_0_0\
        );

    \I__2755\ : InMux
    port map (
            O => \N__14529\,
            I => \N__14523\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14528\,
            I => \N__14511\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14527\,
            I => \N__14507\
        );

    \I__2752\ : InMux
    port map (
            O => \N__14526\,
            I => \N__14504\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__14523\,
            I => \N__14501\
        );

    \I__2750\ : InMux
    port map (
            O => \N__14522\,
            I => \N__14498\
        );

    \I__2749\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14493\
        );

    \I__2748\ : InMux
    port map (
            O => \N__14520\,
            I => \N__14493\
        );

    \I__2747\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14486\
        );

    \I__2746\ : InMux
    port map (
            O => \N__14518\,
            I => \N__14486\
        );

    \I__2745\ : InMux
    port map (
            O => \N__14517\,
            I => \N__14486\
        );

    \I__2744\ : InMux
    port map (
            O => \N__14516\,
            I => \N__14483\
        );

    \I__2743\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14479\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14514\,
            I => \N__14476\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__14511\,
            I => \N__14471\
        );

    \I__2740\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14465\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__14507\,
            I => \N__14460\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__14504\,
            I => \N__14460\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__14501\,
            I => \N__14455\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14498\,
            I => \N__14455\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__14493\,
            I => \N__14450\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__14486\,
            I => \N__14450\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__14483\,
            I => \N__14447\
        );

    \I__2732\ : InMux
    port map (
            O => \N__14482\,
            I => \N__14444\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__14479\,
            I => \N__14441\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__14476\,
            I => \N__14438\
        );

    \I__2729\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14433\
        );

    \I__2728\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14433\
        );

    \I__2727\ : Span4Mux_h
    port map (
            O => \N__14471\,
            I => \N__14430\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14470\,
            I => \N__14425\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14469\,
            I => \N__14425\
        );

    \I__2724\ : InMux
    port map (
            O => \N__14468\,
            I => \N__14422\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14465\,
            I => \N__14419\
        );

    \I__2722\ : Span4Mux_v
    port map (
            O => \N__14460\,
            I => \N__14412\
        );

    \I__2721\ : Span4Mux_h
    port map (
            O => \N__14455\,
            I => \N__14412\
        );

    \I__2720\ : Span4Mux_h
    port map (
            O => \N__14450\,
            I => \N__14412\
        );

    \I__2719\ : Span4Mux_h
    port map (
            O => \N__14447\,
            I => \N__14407\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__14444\,
            I => \N__14407\
        );

    \I__2717\ : Span4Mux_h
    port map (
            O => \N__14441\,
            I => \N__14400\
        );

    \I__2716\ : Span4Mux_v
    port map (
            O => \N__14438\,
            I => \N__14400\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__14433\,
            I => \N__14400\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__14430\,
            I => bu_rx_data_7
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__14425\,
            I => bu_rx_data_7
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__14422\,
            I => bu_rx_data_7
        );

    \I__2711\ : Odrv12
    port map (
            O => \N__14419\,
            I => bu_rx_data_7
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__14412\,
            I => bu_rx_data_7
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__14407\,
            I => bu_rx_data_7
        );

    \I__2708\ : Odrv4
    port map (
            O => \N__14400\,
            I => bu_rx_data_7
        );

    \I__2707\ : InMux
    port map (
            O => \N__14385\,
            I => \N__14375\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14384\,
            I => \N__14375\
        );

    \I__2705\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14367\
        );

    \I__2704\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14361\
        );

    \I__2703\ : InMux
    port map (
            O => \N__14381\,
            I => \N__14361\
        );

    \I__2702\ : InMux
    port map (
            O => \N__14380\,
            I => \N__14358\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__14375\,
            I => \N__14355\
        );

    \I__2700\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14348\
        );

    \I__2699\ : InMux
    port map (
            O => \N__14373\,
            I => \N__14348\
        );

    \I__2698\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14348\
        );

    \I__2697\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14345\
        );

    \I__2696\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14342\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__14367\,
            I => \N__14339\
        );

    \I__2694\ : InMux
    port map (
            O => \N__14366\,
            I => \N__14335\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__14361\,
            I => \N__14332\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__14358\,
            I => \N__14323\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__14355\,
            I => \N__14323\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__14348\,
            I => \N__14323\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__14345\,
            I => \N__14323\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__14342\,
            I => \N__14320\
        );

    \I__2687\ : Span4Mux_v
    port map (
            O => \N__14339\,
            I => \N__14317\
        );

    \I__2686\ : InMux
    port map (
            O => \N__14338\,
            I => \N__14314\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__14335\,
            I => \N__14311\
        );

    \I__2684\ : Span4Mux_v
    port map (
            O => \N__14332\,
            I => \N__14306\
        );

    \I__2683\ : Span4Mux_h
    port map (
            O => \N__14323\,
            I => \N__14306\
        );

    \I__2682\ : Span4Mux_h
    port map (
            O => \N__14320\,
            I => \N__14299\
        );

    \I__2681\ : Span4Mux_h
    port map (
            O => \N__14317\,
            I => \N__14299\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__14314\,
            I => \N__14299\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__14311\,
            I => \N_232\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__14306\,
            I => \N_232\
        );

    \I__2677\ : Odrv4
    port map (
            O => \N__14299\,
            I => \N_232\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14292\,
            I => \N__14289\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__14289\,
            I => \N__14286\
        );

    \I__2674\ : Span4Mux_v
    port map (
            O => \N__14286\,
            I => \N__14283\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__14283\,
            I => \Lab_UT.scctrl.g0_2_0\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__14280\,
            I => \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_1_3_cascade_\
        );

    \I__2671\ : InMux
    port map (
            O => \N__14277\,
            I => \N__14274\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__14274\,
            I => \N__14271\
        );

    \I__2669\ : Odrv12
    port map (
            O => \N__14271\,
            I => \Lab_UT.scctrl.next_state_0_0\
        );

    \I__2668\ : InMux
    port map (
            O => \N__14268\,
            I => \N__14265\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__14265\,
            I => \Lab_UT.scctrl.g0_1_i_0\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__14262\,
            I => \Lab_UT.scctrl.g0_1_i_2_cascade_\
        );

    \I__2665\ : InMux
    port map (
            O => \N__14259\,
            I => \N__14256\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__14256\,
            I => \Lab_UT.scctrl.g0_1_i_4\
        );

    \I__2663\ : InMux
    port map (
            O => \N__14253\,
            I => \N__14250\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__14250\,
            I => \N__14247\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__14247\,
            I => \Lab_UT.scctrl.next_state_rst_2_0\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__14244\,
            I => \Lab_UT.scctrl.G_24_i_a3_0_cascade_\
        );

    \I__2659\ : InMux
    port map (
            O => \N__14241\,
            I => \N__14238\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__14238\,
            I => \Lab_UT.scctrl.N_8\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__14235\,
            I => \Lab_UT.scctrl.N_290_2_cascade_\
        );

    \I__2656\ : InMux
    port map (
            O => \N__14232\,
            I => \N__14229\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__14229\,
            I => \Lab_UT.scctrl.N_8_3\
        );

    \I__2654\ : InMux
    port map (
            O => \N__14226\,
            I => \N__14223\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__14223\,
            I => \Lab_UT.scctrl.g0_1_2_0\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__14220\,
            I => \Lab_UT.scctrl.g3_cascade_\
        );

    \I__2651\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14214\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__14214\,
            I => \Lab_UT.scctrl.g0_1_4\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__14211\,
            I => \Lab_UT.scctrl.next_state_rst_1_cascade_\
        );

    \I__2648\ : InMux
    port map (
            O => \N__14208\,
            I => \N__14205\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__14205\,
            I => \N__14202\
        );

    \I__2646\ : Span4Mux_v
    port map (
            O => \N__14202\,
            I => \N__14199\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__14199\,
            I => \Lab_UT.scctrl.g0_i_0\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__14196\,
            I => \N__14193\
        );

    \I__2643\ : InMux
    port map (
            O => \N__14193\,
            I => \N__14190\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__14190\,
            I => \N__14187\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__14187\,
            I => \Lab_UT.scctrl.g3_0\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__14184\,
            I => \Lab_UT.scctrl.next_state_rst_0_7_cascade_\
        );

    \I__2639\ : InMux
    port map (
            O => \N__14181\,
            I => \N__14178\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__14178\,
            I => \Lab_UT.scctrl.N_10\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__14175\,
            I => \Lab_UT.scctrl.g1_0_4_cascade_\
        );

    \I__2636\ : InMux
    port map (
            O => \N__14172\,
            I => \N__14169\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__14169\,
            I => \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_3\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__14166\,
            I => \Lab_UT.scctrl.N_290_cascade_\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__14163\,
            I => \Lab_UT.scctrl.N_9_cascade_\
        );

    \I__2632\ : InMux
    port map (
            O => \N__14160\,
            I => \N__14157\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__14157\,
            I => \Lab_UT.scctrl.g0_9_0\
        );

    \I__2630\ : InMux
    port map (
            O => \N__14154\,
            I => \N__14151\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__14151\,
            I => \N__14147\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__14150\,
            I => \N__14144\
        );

    \I__2627\ : Span12Mux_v
    port map (
            O => \N__14147\,
            I => \N__14141\
        );

    \I__2626\ : InMux
    port map (
            O => \N__14144\,
            I => \N__14138\
        );

    \I__2625\ : Odrv12
    port map (
            O => \N__14141\,
            I => \Lab_UT.scdp.key1_7\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__14138\,
            I => \Lab_UT.scdp.key1_7\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__14133\,
            I => \N__14129\
        );

    \I__2622\ : InMux
    port map (
            O => \N__14132\,
            I => \N__14126\
        );

    \I__2621\ : InMux
    port map (
            O => \N__14129\,
            I => \N__14123\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__14126\,
            I => \Lab_UT.scdp.key1_0\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__14123\,
            I => \Lab_UT.scdp.key1_0\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__14118\,
            I => \N__14114\
        );

    \I__2617\ : InMux
    port map (
            O => \N__14117\,
            I => \N__14111\
        );

    \I__2616\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14108\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__14111\,
            I => \Lab_UT.scdp.key1_3\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__14108\,
            I => \Lab_UT.scdp.key1_3\
        );

    \I__2613\ : InMux
    port map (
            O => \N__14103\,
            I => \N__14100\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__14100\,
            I => \N__14096\
        );

    \I__2611\ : InMux
    port map (
            O => \N__14099\,
            I => \N__14093\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__14096\,
            I => \Lab_UT.scdp.key2_6\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__14093\,
            I => \Lab_UT.scdp.key2_6\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__14088\,
            I => \N__14084\
        );

    \I__2607\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14081\
        );

    \I__2606\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14078\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__14081\,
            I => \Lab_UT.scdp.key2_4\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__14078\,
            I => \Lab_UT.scdp.key2_4\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__14073\,
            I => \N__14069\
        );

    \I__2602\ : InMux
    port map (
            O => \N__14072\,
            I => \N__14066\
        );

    \I__2601\ : InMux
    port map (
            O => \N__14069\,
            I => \N__14063\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__14066\,
            I => \Lab_UT.scdp.key2_2\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__14063\,
            I => \Lab_UT.scdp.key2_2\
        );

    \I__2598\ : InMux
    port map (
            O => \N__14058\,
            I => \N__14055\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__14055\,
            I => \N__14052\
        );

    \I__2596\ : Span4Mux_s2_v
    port map (
            O => \N__14052\,
            I => \N__14048\
        );

    \I__2595\ : InMux
    port map (
            O => \N__14051\,
            I => \N__14045\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__14048\,
            I => \Lab_UT.scdp.key1_2\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__14045\,
            I => \Lab_UT.scdp.key1_2\
        );

    \I__2592\ : InMux
    port map (
            O => \N__14040\,
            I => \N__14037\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__14037\,
            I => \N__14033\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__14036\,
            I => \N__14030\
        );

    \I__2589\ : Span4Mux_h
    port map (
            O => \N__14033\,
            I => \N__14027\
        );

    \I__2588\ : InMux
    port map (
            O => \N__14030\,
            I => \N__14024\
        );

    \I__2587\ : Odrv4
    port map (
            O => \N__14027\,
            I => \Lab_UT.scdp.key2_5\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__14024\,
            I => \Lab_UT.scdp.key2_5\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__14019\,
            I => \N__14015\
        );

    \I__2584\ : InMux
    port map (
            O => \N__14018\,
            I => \N__14012\
        );

    \I__2583\ : InMux
    port map (
            O => \N__14015\,
            I => \N__14009\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__14012\,
            I => \Lab_UT.scdp.key1_4\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__14009\,
            I => \Lab_UT.scdp.key1_4\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__14004\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_cascade_\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__14001\,
            I => \N__13997\
        );

    \I__2578\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13994\
        );

    \I__2577\ : InMux
    port map (
            O => \N__13997\,
            I => \N__13991\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__13994\,
            I => \N__13988\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__13991\,
            I => \N__13985\
        );

    \I__2574\ : Span4Mux_h
    port map (
            O => \N__13988\,
            I => \N__13981\
        );

    \I__2573\ : Span4Mux_v
    port map (
            O => \N__13985\,
            I => \N__13978\
        );

    \I__2572\ : InMux
    port map (
            O => \N__13984\,
            I => \N__13975\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__13981\,
            I => \Lab_UT.scctrl.N_351\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__13978\,
            I => \Lab_UT.scctrl.N_351\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__13975\,
            I => \Lab_UT.scctrl.N_351\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13968\,
            I => \N__13965\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__13965\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__13962\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_0_0_cascade_\
        );

    \I__2565\ : InMux
    port map (
            O => \N__13959\,
            I => \N__13956\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__13956\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_2\
        );

    \I__2563\ : InMux
    port map (
            O => \N__13953\,
            I => \N__13950\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__13950\,
            I => \N__13947\
        );

    \I__2561\ : Odrv12
    port map (
            O => \N__13947\,
            I => \Lab_UT.scctrl.N_6_2\
        );

    \I__2560\ : InMux
    port map (
            O => \N__13944\,
            I => \N__13941\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__13941\,
            I => \Lab_UT.scctrl.g0_8_1_0\
        );

    \I__2558\ : InMux
    port map (
            O => \N__13938\,
            I => \N__13935\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__13935\,
            I => \N__13932\
        );

    \I__2556\ : Odrv4
    port map (
            O => \N__13932\,
            I => \Lab_UT.scctrl.N_404_2\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__13929\,
            I => \Lab_UT.scctrl.g0_8_1_cascade_\
        );

    \I__2554\ : InMux
    port map (
            O => \N__13926\,
            I => \N__13922\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__13925\,
            I => \N__13919\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__13922\,
            I => \N__13916\
        );

    \I__2551\ : InMux
    port map (
            O => \N__13919\,
            I => \N__13913\
        );

    \I__2550\ : Odrv12
    port map (
            O => \N__13916\,
            I => \Lab_UT.scdp.key1_6\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__13913\,
            I => \Lab_UT.scdp.key1_6\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__13908\,
            I => \Lab_UT.N_100_i_cascade_\
        );

    \I__2547\ : CEMux
    port map (
            O => \N__13905\,
            I => \N__13902\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__13902\,
            I => \N__13899\
        );

    \I__2545\ : Odrv12
    port map (
            O => \N__13899\,
            I => \Lab_UT.scdp.u2.N_100_i_0\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__13896\,
            I => \Lab_UT.scctrl.N_13_0_cascade_\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__13893\,
            I => \Lab_UT.scctrl.N_404_3_cascade_\
        );

    \I__2542\ : InMux
    port map (
            O => \N__13890\,
            I => \N__13877\
        );

    \I__2541\ : InMux
    port map (
            O => \N__13889\,
            I => \N__13877\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13888\,
            I => \N__13877\
        );

    \I__2539\ : InMux
    port map (
            O => \N__13887\,
            I => \N__13877\
        );

    \I__2538\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13874\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__13877\,
            I => \buart.Z_rx.N_80\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__13874\,
            I => \buart.Z_rx.N_80\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13869\,
            I => \N__13866\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__13866\,
            I => \N__13862\
        );

    \I__2533\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13854\
        );

    \I__2532\ : Span4Mux_h
    port map (
            O => \N__13862\,
            I => \N__13851\
        );

    \I__2531\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13848\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13860\,
            I => \N__13843\
        );

    \I__2529\ : InMux
    port map (
            O => \N__13859\,
            I => \N__13843\
        );

    \I__2528\ : InMux
    port map (
            O => \N__13858\,
            I => \N__13838\
        );

    \I__2527\ : InMux
    port map (
            O => \N__13857\,
            I => \N__13838\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13854\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__13851\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__13848\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__13843\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__13838\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__13827\,
            I => \N__13823\
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__13826\,
            I => \N__13817\
        );

    \I__2519\ : InMux
    port map (
            O => \N__13823\,
            I => \N__13814\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13822\,
            I => \N__13811\
        );

    \I__2517\ : InMux
    port map (
            O => \N__13821\,
            I => \N__13808\
        );

    \I__2516\ : InMux
    port map (
            O => \N__13820\,
            I => \N__13803\
        );

    \I__2515\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13803\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__13814\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__13811\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__13808\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__13803\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13794\,
            I => \N__13787\
        );

    \I__2509\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13784\
        );

    \I__2508\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13781\
        );

    \I__2507\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13776\
        );

    \I__2506\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13776\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13787\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__13784\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__13781\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__13776\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13767\,
            I => \N__13757\
        );

    \I__2500\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13757\
        );

    \I__2499\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13757\
        );

    \I__2498\ : InMux
    port map (
            O => \N__13764\,
            I => \N__13754\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__13757\,
            I => \buart__rx_N_86_i_0_o2_1_0\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__13754\,
            I => \buart__rx_N_86_i_0_o2_1_0\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13744\
        );

    \I__2494\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13739\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13739\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__13744\,
            I => \N__13736\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__13739\,
            I => \Lab_UT.N_252\
        );

    \I__2490\ : Odrv4
    port map (
            O => \N__13736\,
            I => \Lab_UT.N_252\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__13731\,
            I => \N__13727\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__13730\,
            I => \N__13718\
        );

    \I__2487\ : InMux
    port map (
            O => \N__13727\,
            I => \N__13713\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13726\,
            I => \N__13710\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13703\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13703\
        );

    \I__2483\ : InMux
    port map (
            O => \N__13723\,
            I => \N__13703\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13694\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13694\
        );

    \I__2480\ : InMux
    port map (
            O => \N__13718\,
            I => \N__13694\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13717\,
            I => \N__13694\
        );

    \I__2478\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13691\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__13713\,
            I => \buart__rx_bitcount_4\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__13710\,
            I => \buart__rx_bitcount_4\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__13703\,
            I => \buart__rx_bitcount_4\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__13694\,
            I => \buart__rx_bitcount_4\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__13691\,
            I => \buart__rx_bitcount_4\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__13680\,
            I => \buart__rx_N_86_i_0_o2_1_0_cascade_\
        );

    \I__2471\ : InMux
    port map (
            O => \N__13677\,
            I => \N__13664\
        );

    \I__2470\ : InMux
    port map (
            O => \N__13676\,
            I => \N__13661\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13658\
        );

    \I__2468\ : InMux
    port map (
            O => \N__13674\,
            I => \N__13649\
        );

    \I__2467\ : InMux
    port map (
            O => \N__13673\,
            I => \N__13649\
        );

    \I__2466\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13649\
        );

    \I__2465\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13649\
        );

    \I__2464\ : InMux
    port map (
            O => \N__13670\,
            I => \N__13646\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13669\,
            I => \N__13639\
        );

    \I__2462\ : InMux
    port map (
            O => \N__13668\,
            I => \N__13639\
        );

    \I__2461\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13639\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__13664\,
            I => \buart__rx_bitcount_1\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__13661\,
            I => \buart__rx_bitcount_1\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__13658\,
            I => \buart__rx_bitcount_1\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__13649\,
            I => \buart__rx_bitcount_1\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__13646\,
            I => \buart__rx_bitcount_1\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__13639\,
            I => \buart__rx_bitcount_1\
        );

    \I__2454\ : InMux
    port map (
            O => \N__13626\,
            I => \N__13623\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__13623\,
            I => \N__13620\
        );

    \I__2452\ : Span4Mux_h
    port map (
            O => \N__13620\,
            I => \N__13617\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__13617\,
            I => \Lab_UT.scctrl.r4.delay4\
        );

    \I__2450\ : InMux
    port map (
            O => \N__13614\,
            I => \N__13611\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13611\,
            I => \N__13607\
        );

    \I__2448\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13604\
        );

    \I__2447\ : Span4Mux_h
    port map (
            O => \N__13607\,
            I => \N__13601\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__13604\,
            I => \Lab_UT.scctrl.delay3\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__13601\,
            I => \Lab_UT.scctrl.delay3\
        );

    \I__2444\ : InMux
    port map (
            O => \N__13596\,
            I => \N__13593\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__13593\,
            I => \Lab_UT.scctrl.delay1\
        );

    \I__2442\ : InMux
    port map (
            O => \N__13590\,
            I => \N__13587\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__13587\,
            I => \Lab_UT.scctrl.delay2\
        );

    \I__2440\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13581\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__13581\,
            I => \Lab_UT.scctrl.N_384\
        );

    \I__2438\ : InMux
    port map (
            O => \N__13578\,
            I => \N__13572\
        );

    \I__2437\ : InMux
    port map (
            O => \N__13577\,
            I => \N__13572\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__13572\,
            I => \N__13569\
        );

    \I__2435\ : Odrv12
    port map (
            O => \N__13569\,
            I => \Lab_UT.scctrl.N_385\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__13566\,
            I => \Lab_UT.scctrl.N_384_cascade_\
        );

    \I__2433\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13559\
        );

    \I__2432\ : InMux
    port map (
            O => \N__13562\,
            I => \N__13556\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__13559\,
            I => \buart__rx_shifter_0_fast_2\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__13556\,
            I => \buart__rx_shifter_0_fast_2\
        );

    \I__2429\ : InMux
    port map (
            O => \N__13551\,
            I => \N__13542\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__13550\,
            I => \N__13538\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__13549\,
            I => \N__13534\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13548\,
            I => \N__13531\
        );

    \I__2425\ : InMux
    port map (
            O => \N__13547\,
            I => \N__13524\
        );

    \I__2424\ : InMux
    port map (
            O => \N__13546\,
            I => \N__13524\
        );

    \I__2423\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13524\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__13542\,
            I => \N__13521\
        );

    \I__2421\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13518\
        );

    \I__2420\ : InMux
    port map (
            O => \N__13538\,
            I => \N__13510\
        );

    \I__2419\ : InMux
    port map (
            O => \N__13537\,
            I => \N__13510\
        );

    \I__2418\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13510\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__13531\,
            I => \N__13505\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__13524\,
            I => \N__13502\
        );

    \I__2415\ : Span4Mux_v
    port map (
            O => \N__13521\,
            I => \N__13498\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__13518\,
            I => \N__13495\
        );

    \I__2413\ : CascadeMux
    port map (
            O => \N__13517\,
            I => \N__13491\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__13510\,
            I => \N__13488\
        );

    \I__2411\ : InMux
    port map (
            O => \N__13509\,
            I => \N__13483\
        );

    \I__2410\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13483\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__13505\,
            I => \N__13478\
        );

    \I__2408\ : Span4Mux_v
    port map (
            O => \N__13502\,
            I => \N__13478\
        );

    \I__2407\ : InMux
    port map (
            O => \N__13501\,
            I => \N__13475\
        );

    \I__2406\ : Span4Mux_h
    port map (
            O => \N__13498\,
            I => \N__13470\
        );

    \I__2405\ : Span4Mux_v
    port map (
            O => \N__13495\,
            I => \N__13470\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13494\,
            I => \N__13465\
        );

    \I__2403\ : InMux
    port map (
            O => \N__13491\,
            I => \N__13465\
        );

    \I__2402\ : Span4Mux_s2_v
    port map (
            O => \N__13488\,
            I => \N__13462\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__13483\,
            I => bu_rx_data_3
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__13478\,
            I => bu_rx_data_3
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__13475\,
            I => bu_rx_data_3
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__13470\,
            I => bu_rx_data_3
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__13465\,
            I => bu_rx_data_3
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__13462\,
            I => bu_rx_data_3
        );

    \I__2395\ : CEMux
    port map (
            O => \N__13449\,
            I => \N__13422\
        );

    \I__2394\ : CEMux
    port map (
            O => \N__13448\,
            I => \N__13422\
        );

    \I__2393\ : CEMux
    port map (
            O => \N__13447\,
            I => \N__13422\
        );

    \I__2392\ : CEMux
    port map (
            O => \N__13446\,
            I => \N__13422\
        );

    \I__2391\ : CEMux
    port map (
            O => \N__13445\,
            I => \N__13422\
        );

    \I__2390\ : CEMux
    port map (
            O => \N__13444\,
            I => \N__13422\
        );

    \I__2389\ : CEMux
    port map (
            O => \N__13443\,
            I => \N__13422\
        );

    \I__2388\ : CEMux
    port map (
            O => \N__13442\,
            I => \N__13422\
        );

    \I__2387\ : CEMux
    port map (
            O => \N__13441\,
            I => \N__13422\
        );

    \I__2386\ : GlobalMux
    port map (
            O => \N__13422\,
            I => \N__13419\
        );

    \I__2385\ : gio2CtrlBuf
    port map (
            O => \N__13419\,
            I => \N_76_i_g\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__13416\,
            I => \buart.Z_rx.bitcountN11_15_i_0_o2_0_cascade_\
        );

    \I__2383\ : InMux
    port map (
            O => \N__13413\,
            I => \N__13408\
        );

    \I__2382\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13405\
        );

    \I__2381\ : InMux
    port map (
            O => \N__13411\,
            I => \N__13401\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__13408\,
            I => \N__13393\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__13405\,
            I => \N__13393\
        );

    \I__2378\ : InMux
    port map (
            O => \N__13404\,
            I => \N__13390\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__13401\,
            I => \N__13387\
        );

    \I__2376\ : InMux
    port map (
            O => \N__13400\,
            I => \N__13384\
        );

    \I__2375\ : InMux
    port map (
            O => \N__13399\,
            I => \N__13379\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13398\,
            I => \N__13379\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__13393\,
            I => \N__13376\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__13390\,
            I => \N__13373\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__13387\,
            I => \Lab_UT.scctrl.N_241\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__13384\,
            I => \Lab_UT.scctrl.N_241\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__13379\,
            I => \Lab_UT.scctrl.N_241\
        );

    \I__2368\ : Odrv4
    port map (
            O => \N__13376\,
            I => \Lab_UT.scctrl.N_241\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__13373\,
            I => \Lab_UT.scctrl.N_241\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__13362\,
            I => \Lab_UT.scctrl.g0_70_1_cascade_\
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__13359\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0_cascade_\
        );

    \I__2364\ : InMux
    port map (
            O => \N__13356\,
            I => \N__13349\
        );

    \I__2363\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13349\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__13354\,
            I => \N__13346\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__13349\,
            I => \N__13342\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13346\,
            I => \N__13337\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13345\,
            I => \N__13337\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__13342\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__13337\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0\
        );

    \I__2356\ : InMux
    port map (
            O => \N__13332\,
            I => \N__13329\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__13329\,
            I => \buart__rx_shifter_2_fast_6\
        );

    \I__2354\ : InMux
    port map (
            O => \N__13326\,
            I => \N__13317\
        );

    \I__2353\ : InMux
    port map (
            O => \N__13325\,
            I => \N__13317\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13324\,
            I => \N__13317\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__13317\,
            I => \Lab_UT.scctrl.N_444\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__13314\,
            I => \N__13310\
        );

    \I__2349\ : InMux
    port map (
            O => \N__13313\,
            I => \N__13305\
        );

    \I__2348\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13305\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__13305\,
            I => bu_rx_data_i_2_fast_3
        );

    \I__2346\ : InMux
    port map (
            O => \N__13302\,
            I => \N__13299\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__13299\,
            I => \N__13296\
        );

    \I__2344\ : Span4Mux_h
    port map (
            O => \N__13296\,
            I => \N__13293\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__13293\,
            I => \N_243_reti\
        );

    \I__2342\ : InMux
    port map (
            O => \N__13290\,
            I => \N__13287\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__13287\,
            I => \Lab_UT.scctrl.N_219i\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__13284\,
            I => \N__13281\
        );

    \I__2339\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13278\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__13278\,
            I => \Lab_UT.scctrl.N_271_0_0\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__13275\,
            I => \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_1_cascade_\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13272\,
            I => \N__13269\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__13269\,
            I => \Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__13266\,
            I => \Lab_UT.scctrl.g0_i_o7_1_cascade_\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__13263\,
            I => \Lab_UT.scctrl.N_12_2_cascade_\
        );

    \I__2332\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13255\
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__13259\,
            I => \N__13251\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13247\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13255\,
            I => \N__13244\
        );

    \I__2328\ : InMux
    port map (
            O => \N__13254\,
            I => \N__13241\
        );

    \I__2327\ : InMux
    port map (
            O => \N__13251\,
            I => \N__13238\
        );

    \I__2326\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13235\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__13247\,
            I => bu_rx_data_i_2_3_rep1
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__13244\,
            I => bu_rx_data_i_2_3_rep1
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__13241\,
            I => bu_rx_data_i_2_3_rep1
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__13238\,
            I => bu_rx_data_i_2_3_rep1
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__13235\,
            I => bu_rx_data_i_2_3_rep1
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__13224\,
            I => \N__13220\
        );

    \I__2319\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13216\
        );

    \I__2318\ : InMux
    port map (
            O => \N__13220\,
            I => \N__13211\
        );

    \I__2317\ : InMux
    port map (
            O => \N__13219\,
            I => \N__13211\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__13216\,
            I => \N__13208\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__13211\,
            I => \N__13205\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__13208\,
            I => \Lab_UT.scctrl.N_259\
        );

    \I__2313\ : Odrv12
    port map (
            O => \N__13205\,
            I => \Lab_UT.scctrl.N_259\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__13200\,
            I => \N__13197\
        );

    \I__2311\ : InMux
    port map (
            O => \N__13197\,
            I => \N__13194\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__13194\,
            I => \N__13191\
        );

    \I__2309\ : Span4Mux_h
    port map (
            O => \N__13191\,
            I => \N__13188\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__13188\,
            I => \Lab_UT.scctrl.g0_1_i_a8_0_1\
        );

    \I__2307\ : InMux
    port map (
            O => \N__13185\,
            I => \N__13182\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__13182\,
            I => \Lab_UT.scctrl.N_7_0\
        );

    \I__2305\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13176\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__13176\,
            I => \Lab_UT.scctrl.N_10_0\
        );

    \I__2303\ : InMux
    port map (
            O => \N__13173\,
            I => \N__13165\
        );

    \I__2302\ : InMux
    port map (
            O => \N__13172\,
            I => \N__13165\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13171\,
            I => \N__13162\
        );

    \I__2300\ : InMux
    port map (
            O => \N__13170\,
            I => \N__13159\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__13165\,
            I => \N__13156\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__13162\,
            I => \Lab_UT.scctrl.N_219\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__13159\,
            I => \Lab_UT.scctrl.N_219\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__13156\,
            I => \Lab_UT.scctrl.N_219\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__13149\,
            I => \N__13145\
        );

    \I__2294\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13139\
        );

    \I__2293\ : InMux
    port map (
            O => \N__13145\,
            I => \N__13139\
        );

    \I__2292\ : InMux
    port map (
            O => \N__13144\,
            I => \N__13136\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__13139\,
            I => \N__13133\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__13136\,
            I => \buart__rx_shifter_0_fast_1\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__13133\,
            I => \buart__rx_shifter_0_fast_1\
        );

    \I__2288\ : InMux
    port map (
            O => \N__13128\,
            I => \N__13125\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__13125\,
            I => \Lab_UT.scctrl.g0_0_i_0\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__13122\,
            I => \Lab_UT.scctrl.g0_0_i_1_cascade_\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__13119\,
            I => \Lab_UT.scctrl.g0_0_i_1_0_cascade_\
        );

    \I__2284\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13113\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__13113\,
            I => \Lab_UT.scctrl.N_5_1\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__13110\,
            I => \Lab_UT.scctrl.g0_2_0_0_a3_1_1_cascade_\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__13107\,
            I => \Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0_cascade_\
        );

    \I__2280\ : InMux
    port map (
            O => \N__13104\,
            I => \N__13101\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__13101\,
            I => \Lab_UT.scctrl.g1_0_5\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__13098\,
            I => \Lab_UT.scctrl.next_state_1_0_2_cascade_\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__13095\,
            I => \Lab_UT.scctrl.N_444_0_cascade_\
        );

    \I__2276\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13089\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__13089\,
            I => \Lab_UT.scctrl.N_319_1_0\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__13086\,
            I => \Lab_UT.scctrl.N_223_1_0_cascade_\
        );

    \I__2273\ : InMux
    port map (
            O => \N__13083\,
            I => \N__13080\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__13080\,
            I => \Lab_UT.scctrl.N_414_1_0\
        );

    \I__2271\ : InMux
    port map (
            O => \N__13077\,
            I => \N__13074\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__13074\,
            I => \Lab_UT.scctrl.N_444_0\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__13071\,
            I => \Lab_UT.scctrl.N_223_1_cascade_\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__13068\,
            I => \Lab_UT.scctrl.N_414_1_cascade_\
        );

    \I__2267\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13062\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__13062\,
            I => \N__13058\
        );

    \I__2265\ : InMux
    port map (
            O => \N__13061\,
            I => \N__13055\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__13058\,
            I => \Lab_UT.scctrl.g1_0_2_0\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__13055\,
            I => \Lab_UT.scctrl.g1_0_2_0\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__13050\,
            I => \Lab_UT.scctrl.next_state_1_2_cascade_\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__13047\,
            I => \Lab_UT.scctrl.N_534_reti_cascade_\
        );

    \I__2260\ : InMux
    port map (
            O => \N__13044\,
            I => \N__13041\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__13041\,
            I => \Lab_UT.scctrl.N_266i\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__13038\,
            I => \N__13034\
        );

    \I__2257\ : InMux
    port map (
            O => \N__13037\,
            I => \N__13027\
        );

    \I__2256\ : InMux
    port map (
            O => \N__13034\,
            I => \N__13024\
        );

    \I__2255\ : InMux
    port map (
            O => \N__13033\,
            I => \N__13021\
        );

    \I__2254\ : InMux
    port map (
            O => \N__13032\,
            I => \N__13014\
        );

    \I__2253\ : InMux
    port map (
            O => \N__13031\,
            I => \N__13011\
        );

    \I__2252\ : InMux
    port map (
            O => \N__13030\,
            I => \N__13007\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__13027\,
            I => \N__13004\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__13024\,
            I => \N__13001\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__13021\,
            I => \N__12998\
        );

    \I__2248\ : InMux
    port map (
            O => \N__13020\,
            I => \N__12993\
        );

    \I__2247\ : InMux
    port map (
            O => \N__13019\,
            I => \N__12993\
        );

    \I__2246\ : InMux
    port map (
            O => \N__13018\,
            I => \N__12988\
        );

    \I__2245\ : InMux
    port map (
            O => \N__13017\,
            I => \N__12988\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__13014\,
            I => \N__12985\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__13011\,
            I => \N__12980\
        );

    \I__2242\ : InMux
    port map (
            O => \N__13010\,
            I => \N__12977\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__13007\,
            I => \N__12971\
        );

    \I__2240\ : Span12Mux_s7_h
    port map (
            O => \N__13004\,
            I => \N__12968\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__13001\,
            I => \N__12957\
        );

    \I__2238\ : Span4Mux_h
    port map (
            O => \N__12998\,
            I => \N__12957\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__12993\,
            I => \N__12957\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__12988\,
            I => \N__12957\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__12985\,
            I => \N__12957\
        );

    \I__2234\ : InMux
    port map (
            O => \N__12984\,
            I => \N__12954\
        );

    \I__2233\ : InMux
    port map (
            O => \N__12983\,
            I => \N__12951\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__12980\,
            I => \N__12946\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__12977\,
            I => \N__12946\
        );

    \I__2230\ : InMux
    port map (
            O => \N__12976\,
            I => \N__12939\
        );

    \I__2229\ : InMux
    port map (
            O => \N__12975\,
            I => \N__12939\
        );

    \I__2228\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12939\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__12971\,
            I => bu_rx_data_2
        );

    \I__2226\ : Odrv12
    port map (
            O => \N__12968\,
            I => bu_rx_data_2
        );

    \I__2225\ : Odrv4
    port map (
            O => \N__12957\,
            I => bu_rx_data_2
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__12954\,
            I => bu_rx_data_2
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__12951\,
            I => bu_rx_data_2
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__12946\,
            I => bu_rx_data_2
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__12939\,
            I => bu_rx_data_2
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__12924\,
            I => \N__12921\
        );

    \I__2219\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12918\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__12918\,
            I => \N__12915\
        );

    \I__2217\ : Span4Mux_v
    port map (
            O => \N__12915\,
            I => \N__12911\
        );

    \I__2216\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12908\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__12911\,
            I => \Lab_UT.N_540\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__12908\,
            I => \Lab_UT.N_540\
        );

    \I__2213\ : InMux
    port map (
            O => \N__12903\,
            I => \N__12900\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__12900\,
            I => \Lab_UT.scctrl.N_399_0\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12897\,
            I => \N__12894\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__12894\,
            I => \Lab_UT.scctrl.sccEldByte_i_a2_0Z0Z_1\
        );

    \I__2209\ : InMux
    port map (
            O => \N__12891\,
            I => \N__12888\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__12888\,
            I => \Lab_UT.scctrl.g2\
        );

    \I__2207\ : InMux
    port map (
            O => \N__12885\,
            I => \N__12882\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__12882\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12875\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__12878\,
            I => \N__12872\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__12875\,
            I => \N__12869\
        );

    \I__2202\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12866\
        );

    \I__2201\ : Odrv4
    port map (
            O => \N__12869\,
            I => \Lab_UT.scdp.key0_4\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__12866\,
            I => \Lab_UT.scdp.key0_4\
        );

    \I__2199\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12855\
        );

    \I__2198\ : InMux
    port map (
            O => \N__12860\,
            I => \N__12855\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__12855\,
            I => \Lab_UT.scdp.prng_lfsr_4\
        );

    \I__2196\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12849\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__12849\,
            I => \N__12845\
        );

    \I__2194\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12842\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__12845\,
            I => \Lab_UT.scdp.key3_4\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__12842\,
            I => \Lab_UT.scdp.key3_4\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12837\,
            I => \N__12834\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__12834\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28\
        );

    \I__2189\ : InMux
    port map (
            O => \N__12831\,
            I => \N__12825\
        );

    \I__2188\ : InMux
    port map (
            O => \N__12830\,
            I => \N__12825\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__12825\,
            I => \N__12822\
        );

    \I__2186\ : Span4Mux_h
    port map (
            O => \N__12822\,
            I => \N__12819\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__12819\,
            I => \Lab_UT.scdp.prng_lfsr_11\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__12816\,
            I => \N__12813\
        );

    \I__2183\ : InMux
    port map (
            O => \N__12813\,
            I => \N__12810\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__12810\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26\
        );

    \I__2181\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12801\
        );

    \I__2180\ : InMux
    port map (
            O => \N__12806\,
            I => \N__12801\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__12801\,
            I => \Lab_UT.scdp.prng_lfsr_12\
        );

    \I__2178\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12795\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__12795\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9\
        );

    \I__2176\ : CEMux
    port map (
            O => \N__12792\,
            I => \N__12765\
        );

    \I__2175\ : CEMux
    port map (
            O => \N__12791\,
            I => \N__12765\
        );

    \I__2174\ : CEMux
    port map (
            O => \N__12790\,
            I => \N__12765\
        );

    \I__2173\ : CEMux
    port map (
            O => \N__12789\,
            I => \N__12765\
        );

    \I__2172\ : CEMux
    port map (
            O => \N__12788\,
            I => \N__12765\
        );

    \I__2171\ : CEMux
    port map (
            O => \N__12787\,
            I => \N__12765\
        );

    \I__2170\ : CEMux
    port map (
            O => \N__12786\,
            I => \N__12765\
        );

    \I__2169\ : CEMux
    port map (
            O => \N__12785\,
            I => \N__12765\
        );

    \I__2168\ : CEMux
    port map (
            O => \N__12784\,
            I => \N__12765\
        );

    \I__2167\ : GlobalMux
    port map (
            O => \N__12765\,
            I => \N__12762\
        );

    \I__2166\ : gio2CtrlBuf
    port map (
            O => \N__12762\,
            I => \Lab_UT.sccLdLFSR_g\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12759\,
            I => \N__12756\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__12756\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__12753\,
            I => \N__12750\
        );

    \I__2162\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12747\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__12747\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24\
        );

    \I__2160\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12741\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__12741\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__12738\,
            I => \Lab_UT.scdp.d2eData_3_0_cascade_\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12735\,
            I => \N__12732\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__12732\,
            I => \N__12729\
        );

    \I__2155\ : Span4Mux_h
    port map (
            O => \N__12729\,
            I => \N__12725\
        );

    \I__2154\ : InMux
    port map (
            O => \N__12728\,
            I => \N__12722\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__12725\,
            I => \Lab_UT.scdp.N_262_i\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__12722\,
            I => \Lab_UT.scdp.N_262_i\
        );

    \I__2151\ : InMux
    port map (
            O => \N__12717\,
            I => \N__12714\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__12714\,
            I => \N__12711\
        );

    \I__2149\ : Odrv12
    port map (
            O => \N__12711\,
            I => \Lab_UT.scdp.u1.g0_0_i_a5_0_0\
        );

    \I__2148\ : InMux
    port map (
            O => \N__12708\,
            I => \N__12702\
        );

    \I__2147\ : InMux
    port map (
            O => \N__12707\,
            I => \N__12702\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__12702\,
            I => \N__12699\
        );

    \I__2145\ : Span4Mux_h
    port map (
            O => \N__12699\,
            I => \N__12695\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12698\,
            I => \N__12692\
        );

    \I__2143\ : Span4Mux_v
    port map (
            O => \N__12695\,
            I => \N__12687\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__12692\,
            I => \N__12684\
        );

    \I__2141\ : InMux
    port map (
            O => \N__12691\,
            I => \N__12679\
        );

    \I__2140\ : InMux
    port map (
            O => \N__12690\,
            I => \N__12679\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__12687\,
            I => \Lab_UT.scdp.d2eData_3_0\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__12684\,
            I => \Lab_UT.scdp.d2eData_3_0\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__12679\,
            I => \Lab_UT.scdp.d2eData_3_0\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__12672\,
            I => \N__12668\
        );

    \I__2135\ : InMux
    port map (
            O => \N__12671\,
            I => \N__12660\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12668\,
            I => \N__12660\
        );

    \I__2133\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12655\
        );

    \I__2132\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12655\
        );

    \I__2131\ : InMux
    port map (
            O => \N__12665\,
            I => \N__12652\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__12660\,
            I => \N__12649\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__12655\,
            I => \N__12646\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__12652\,
            I => \Lab_UT.scdp.u1.byteToDecryptZ0Z_2\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__12649\,
            I => \Lab_UT.scdp.u1.byteToDecryptZ0Z_2\
        );

    \I__2126\ : Odrv12
    port map (
            O => \N__12646\,
            I => \Lab_UT.scdp.u1.byteToDecryptZ0Z_2\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12639\,
            I => \N__12627\
        );

    \I__2124\ : InMux
    port map (
            O => \N__12638\,
            I => \N__12627\
        );

    \I__2123\ : InMux
    port map (
            O => \N__12637\,
            I => \N__12627\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12636\,
            I => \N__12627\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__12627\,
            I => \N__12622\
        );

    \I__2120\ : InMux
    port map (
            O => \N__12626\,
            I => \N__12617\
        );

    \I__2119\ : InMux
    port map (
            O => \N__12625\,
            I => \N__12617\
        );

    \I__2118\ : Span12Mux_s4_h
    port map (
            O => \N__12622\,
            I => \N__12613\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__12617\,
            I => \N__12610\
        );

    \I__2116\ : InMux
    port map (
            O => \N__12616\,
            I => \N__12607\
        );

    \I__2115\ : Odrv12
    port map (
            O => \N__12613\,
            I => \Lab_UT.scdp.d2eData_3_2\
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__12610\,
            I => \Lab_UT.scdp.d2eData_3_2\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__12607\,
            I => \Lab_UT.scdp.d2eData_3_2\
        );

    \I__2112\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12597\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__12597\,
            I => \N__12594\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__12594\,
            I => \Lab_UT.scdp.u1.g0_0_i_a5_0_0_0\
        );

    \I__2109\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12588\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__12588\,
            I => \N__12584\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__12587\,
            I => \N__12581\
        );

    \I__2106\ : Span4Mux_v
    port map (
            O => \N__12584\,
            I => \N__12578\
        );

    \I__2105\ : InMux
    port map (
            O => \N__12581\,
            I => \N__12575\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__12578\,
            I => \Lab_UT.scdp.key0_6\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__12575\,
            I => \Lab_UT.scdp.key0_6\
        );

    \I__2102\ : InMux
    port map (
            O => \N__12570\,
            I => \N__12565\
        );

    \I__2101\ : InMux
    port map (
            O => \N__12569\,
            I => \N__12560\
        );

    \I__2100\ : InMux
    port map (
            O => \N__12568\,
            I => \N__12560\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__12565\,
            I => \N__12557\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__12560\,
            I => \N__12554\
        );

    \I__2097\ : Span4Mux_h
    port map (
            O => \N__12557\,
            I => \N__12551\
        );

    \I__2096\ : Span4Mux_h
    port map (
            O => \N__12554\,
            I => \N__12548\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__12551\,
            I => \Lab_UT.scdp.prng_lfsr_6\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__12548\,
            I => \Lab_UT.scdp.prng_lfsr_6\
        );

    \I__2093\ : InMux
    port map (
            O => \N__12543\,
            I => \N__12540\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__12540\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20\
        );

    \I__2091\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12534\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__12534\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__12531\,
            I => \Lab_UT.scctrl.N_22_i_cascade_\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__12528\,
            I => \Lab_UT.state_1_ret_0_RNI9C1NH_0_cascade_\
        );

    \I__2087\ : InMux
    port map (
            O => \N__12525\,
            I => \N__12521\
        );

    \I__2086\ : InMux
    port map (
            O => \N__12524\,
            I => \N__12518\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__12521\,
            I => \Lab_UT.scdp.key3_5\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__12518\,
            I => \Lab_UT.scdp.key3_5\
        );

    \I__2083\ : InMux
    port map (
            O => \N__12513\,
            I => \N__12504\
        );

    \I__2082\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12504\
        );

    \I__2081\ : InMux
    port map (
            O => \N__12511\,
            I => \N__12504\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__12504\,
            I => \Lab_UT.state_1_ret_0_RNI9C1NH_0\
        );

    \I__2079\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12498\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__12498\,
            I => \N__12494\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__12497\,
            I => \N__12491\
        );

    \I__2076\ : Span4Mux_v
    port map (
            O => \N__12494\,
            I => \N__12488\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12491\,
            I => \N__12485\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__12488\,
            I => \Lab_UT.scdp.key3_6\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__12485\,
            I => \Lab_UT.scdp.key3_6\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12473\
        );

    \I__2071\ : InMux
    port map (
            O => \N__12479\,
            I => \N__12468\
        );

    \I__2070\ : InMux
    port map (
            O => \N__12478\,
            I => \N__12468\
        );

    \I__2069\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12463\
        );

    \I__2068\ : InMux
    port map (
            O => \N__12476\,
            I => \N__12463\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__12473\,
            I => \Lab_UT.state_1_RNI6EDGH_0_2\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__12468\,
            I => \Lab_UT.state_1_RNI6EDGH_0_2\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__12463\,
            I => \Lab_UT.state_1_RNI6EDGH_0_2\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__12456\,
            I => \N__12452\
        );

    \I__2063\ : InMux
    port map (
            O => \N__12455\,
            I => \N__12449\
        );

    \I__2062\ : InMux
    port map (
            O => \N__12452\,
            I => \N__12446\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__12449\,
            I => \Lab_UT.scdp.key0_5\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__12446\,
            I => \Lab_UT.scdp.key0_5\
        );

    \I__2059\ : InMux
    port map (
            O => \N__12441\,
            I => \N__12438\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__12438\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__2057\ : InMux
    port map (
            O => \N__12435\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__2056\ : InMux
    port map (
            O => \N__12432\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__2055\ : CEMux
    port map (
            O => \N__12429\,
            I => \N__12426\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__12426\,
            I => \N__12422\
        );

    \I__2053\ : CEMux
    port map (
            O => \N__12425\,
            I => \N__12419\
        );

    \I__2052\ : Span4Mux_v
    port map (
            O => \N__12422\,
            I => \N__12416\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__12419\,
            I => \N__12413\
        );

    \I__2050\ : Span4Mux_h
    port map (
            O => \N__12416\,
            I => \N__12410\
        );

    \I__2049\ : Sp12to4
    port map (
            O => \N__12413\,
            I => \N__12407\
        );

    \I__2048\ : Odrv4
    port map (
            O => \N__12410\,
            I => \buart.Z_rx.N_78\
        );

    \I__2047\ : Odrv12
    port map (
            O => \N__12407\,
            I => \buart.Z_rx.N_78\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__12402\,
            I => \Lab_UT.scctrl.N_418_0_cascade_\
        );

    \I__2045\ : InMux
    port map (
            O => \N__12399\,
            I => \N__12396\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__12396\,
            I => \Lab_UT.scctrl.g0_2\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__12393\,
            I => \Lab_UT.scctrl.g0_2_cascade_\
        );

    \I__2042\ : InMux
    port map (
            O => \N__12390\,
            I => \N__12384\
        );

    \I__2041\ : InMux
    port map (
            O => \N__12389\,
            I => \N__12384\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__12384\,
            I => \N__12381\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__12381\,
            I => \Lab_UT.scctrl.g1_1\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__12378\,
            I => \Lab_UT.scctrl.N_418_2_0_cascade_\
        );

    \I__2037\ : InMux
    port map (
            O => \N__12375\,
            I => \N__12372\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__12372\,
            I => \N__12369\
        );

    \I__2035\ : Span12Mux_s3_v
    port map (
            O => \N__12369\,
            I => \N__12366\
        );

    \I__2034\ : Odrv12
    port map (
            O => \N__12366\,
            I => \Lab_UT.scctrl.g1_1_2\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__12363\,
            I => \Lab_UT.scctrl.N_39_i_cascade_\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__12360\,
            I => \CONSTANT_ONE_NET_cascade_\
        );

    \I__2031\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12354\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__12354\,
            I => \N__12351\
        );

    \I__2029\ : Span4Mux_v
    port map (
            O => \N__12351\,
            I => \N__12348\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__12348\,
            I => \ufifo.sb_ram512x8_inst_RNIKTQ21\
        );

    \I__2027\ : InMux
    port map (
            O => \N__12345\,
            I => \N__12342\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__12342\,
            I => \N__12339\
        );

    \I__2025\ : Span4Mux_v
    port map (
            O => \N__12339\,
            I => \N__12336\
        );

    \I__2024\ : Span4Mux_h
    port map (
            O => \N__12336\,
            I => \N__12333\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__12333\,
            I => \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1Z0Z_0\
        );

    \I__2022\ : InMux
    port map (
            O => \N__12330\,
            I => \N__12327\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__12327\,
            I => \N__12317\
        );

    \I__2020\ : InMux
    port map (
            O => \N__12326\,
            I => \N__12299\
        );

    \I__2019\ : InMux
    port map (
            O => \N__12325\,
            I => \N__12299\
        );

    \I__2018\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12299\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12299\
        );

    \I__2016\ : InMux
    port map (
            O => \N__12322\,
            I => \N__12299\
        );

    \I__2015\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12294\
        );

    \I__2014\ : InMux
    port map (
            O => \N__12320\,
            I => \N__12294\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__12317\,
            I => \N__12291\
        );

    \I__2012\ : InMux
    port map (
            O => \N__12316\,
            I => \N__12288\
        );

    \I__2011\ : InMux
    port map (
            O => \N__12315\,
            I => \N__12281\
        );

    \I__2010\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12281\
        );

    \I__2009\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12281\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12274\
        );

    \I__2007\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12274\
        );

    \I__2006\ : InMux
    port map (
            O => \N__12310\,
            I => \N__12274\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__12299\,
            I => \N__12269\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__12294\,
            I => \N__12269\
        );

    \I__2003\ : Span4Mux_h
    port map (
            O => \N__12291\,
            I => \N__12264\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__12288\,
            I => \N__12264\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__12281\,
            I => \N_368\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__12274\,
            I => \N_368\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__12269\,
            I => \N_368\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__12264\,
            I => \N_368\
        );

    \I__1997\ : InMux
    port map (
            O => \N__12255\,
            I => \N__12252\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__12252\,
            I => \N__12249\
        );

    \I__1995\ : Span4Mux_h
    port map (
            O => \N__12249\,
            I => \N__12246\
        );

    \I__1994\ : Span4Mux_v
    port map (
            O => \N__12246\,
            I => \N__12243\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__12243\,
            I => utb_txdata_0
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__12240\,
            I => \N__12237\
        );

    \I__1991\ : InMux
    port map (
            O => \N__12237\,
            I => \N__12234\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__12234\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__1989\ : InMux
    port map (
            O => \N__12231\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__12228\,
            I => \N__12225\
        );

    \I__1987\ : InMux
    port map (
            O => \N__12225\,
            I => \N__12222\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__12222\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__1985\ : InMux
    port map (
            O => \N__12219\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__1984\ : InMux
    port map (
            O => \N__12216\,
            I => \N__12213\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__12213\,
            I => \N__12210\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__12210\,
            I => \Lab_UT.scctrl.N_263_0\
        );

    \I__1981\ : InMux
    port map (
            O => \N__12207\,
            I => \N__12204\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__12204\,
            I => \Lab_UT.scctrl.N_233_0\
        );

    \I__1979\ : InMux
    port map (
            O => \N__12201\,
            I => \N__12198\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__12198\,
            I => \Lab_UT.scctrl.N_351_1_0\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__12195\,
            I => \Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_5_1_cascade_\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__12192\,
            I => \N__12189\
        );

    \I__1975\ : InMux
    port map (
            O => \N__12189\,
            I => \N__12185\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__12188\,
            I => \N__12182\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__12185\,
            I => \N__12179\
        );

    \I__1972\ : InMux
    port map (
            O => \N__12182\,
            I => \N__12176\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__12179\,
            I => \Lab_UT.N_540i\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__12176\,
            I => \Lab_UT.N_540i\
        );

    \I__1969\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12168\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__12168\,
            I => \Lab_UT.scctrl.N_266\
        );

    \I__1967\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12161\
        );

    \I__1966\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12158\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__12161\,
            I => \N__12155\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__12158\,
            I => \Lab_UT.scctrl.N_472_0\
        );

    \I__1963\ : Odrv12
    port map (
            O => \N__12155\,
            I => \Lab_UT.scctrl.N_472_0\
        );

    \I__1962\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12147\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__12147\,
            I => \Lab_UT.scctrl.N_241_reti\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__12144\,
            I => \Lab_UT.scctrl.N_241_reti_cascade_\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__12141\,
            I => \N__12138\
        );

    \I__1958\ : InMux
    port map (
            O => \N__12138\,
            I => \N__12135\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__12135\,
            I => \N__12132\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__12132\,
            I => \Lab_UT.scctrl.N_319_0\
        );

    \I__1955\ : InMux
    port map (
            O => \N__12129\,
            I => \N__12126\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__12126\,
            I => \N__12123\
        );

    \I__1953\ : Odrv4
    port map (
            O => \N__12123\,
            I => \Lab_UT.scctrl.N_414_0\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__12120\,
            I => \Lab_UT.scctrl.N_415_1_cascade_\
        );

    \I__1951\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12114\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__12114\,
            I => \Lab_UT.scctrl.g1_0_0_0\
        );

    \I__1949\ : InMux
    port map (
            O => \N__12111\,
            I => \N__12108\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__12108\,
            I => \Lab_UT.scctrl.N_259i\
        );

    \I__1947\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12102\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__12102\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10\
        );

    \I__1945\ : InMux
    port map (
            O => \N__12099\,
            I => \N__12096\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__12096\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__12093\,
            I => \Lab_UT.scdp.d2eData_3_2_cascade_\
        );

    \I__1942\ : InMux
    port map (
            O => \N__12090\,
            I => \N__12085\
        );

    \I__1941\ : InMux
    port map (
            O => \N__12089\,
            I => \N__12082\
        );

    \I__1940\ : InMux
    port map (
            O => \N__12088\,
            I => \N__12078\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__12085\,
            I => \N__12073\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__12082\,
            I => \N__12073\
        );

    \I__1937\ : InMux
    port map (
            O => \N__12081\,
            I => \N__12070\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__12078\,
            I => \N__12067\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__12073\,
            I => \N__12064\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__12070\,
            I => \N__12061\
        );

    \I__1933\ : Span4Mux_v
    port map (
            O => \N__12067\,
            I => \N__12056\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__12064\,
            I => \N__12056\
        );

    \I__1931\ : Span4Mux_h
    port map (
            O => \N__12061\,
            I => \N__12053\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__12056\,
            I => \Lab_UT.scdp.N_234_i\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__12053\,
            I => \Lab_UT.scdp.N_234_i\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__12048\,
            I => \N__12044\
        );

    \I__1927\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12040\
        );

    \I__1926\ : InMux
    port map (
            O => \N__12044\,
            I => \N__12037\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__12043\,
            I => \N__12031\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__12040\,
            I => \N__12026\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__12037\,
            I => \N__12026\
        );

    \I__1922\ : InMux
    port map (
            O => \N__12036\,
            I => \N__12023\
        );

    \I__1921\ : InMux
    port map (
            O => \N__12035\,
            I => \N__12018\
        );

    \I__1920\ : InMux
    port map (
            O => \N__12034\,
            I => \N__12015\
        );

    \I__1919\ : InMux
    port map (
            O => \N__12031\,
            I => \N__12012\
        );

    \I__1918\ : Sp12to4
    port map (
            O => \N__12026\,
            I => \N__12007\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__12023\,
            I => \N__12007\
        );

    \I__1916\ : InMux
    port map (
            O => \N__12022\,
            I => \N__12004\
        );

    \I__1915\ : InMux
    port map (
            O => \N__12021\,
            I => \N__12001\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__12018\,
            I => \Lab_UT.scdp.byteToDecrypt_5\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__12015\,
            I => \Lab_UT.scdp.byteToDecrypt_5\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__12012\,
            I => \Lab_UT.scdp.byteToDecrypt_5\
        );

    \I__1911\ : Odrv12
    port map (
            O => \N__12007\,
            I => \Lab_UT.scdp.byteToDecrypt_5\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__12004\,
            I => \Lab_UT.scdp.byteToDecrypt_5\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__12001\,
            I => \Lab_UT.scdp.byteToDecrypt_5\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11988\,
            I => \N__11985\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__11985\,
            I => \N__11982\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__11982\,
            I => \Lab_UT.scdp.N_228_i_0\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__11979\,
            I => \Lab_UT.scdp.g0_0_i_0_cascade_\
        );

    \I__1904\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11964\
        );

    \I__1903\ : InMux
    port map (
            O => \N__11975\,
            I => \N__11964\
        );

    \I__1902\ : InMux
    port map (
            O => \N__11974\,
            I => \N__11964\
        );

    \I__1901\ : InMux
    port map (
            O => \N__11973\,
            I => \N__11959\
        );

    \I__1900\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11956\
        );

    \I__1899\ : InMux
    port map (
            O => \N__11971\,
            I => \N__11952\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__11964\,
            I => \N__11949\
        );

    \I__1897\ : InMux
    port map (
            O => \N__11963\,
            I => \N__11946\
        );

    \I__1896\ : InMux
    port map (
            O => \N__11962\,
            I => \N__11943\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__11959\,
            I => \N__11938\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__11956\,
            I => \N__11938\
        );

    \I__1893\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11935\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__11952\,
            I => \Lab_UT.scdp.d2eData_3_5\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__11949\,
            I => \Lab_UT.scdp.d2eData_3_5\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__11946\,
            I => \Lab_UT.scdp.d2eData_3_5\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__11943\,
            I => \Lab_UT.scdp.d2eData_3_5\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__11938\,
            I => \Lab_UT.scdp.d2eData_3_5\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__11935\,
            I => \Lab_UT.scdp.d2eData_3_5\
        );

    \I__1886\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11919\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__11919\,
            I => \N__11916\
        );

    \I__1884\ : Span4Mux_h
    port map (
            O => \N__11916\,
            I => \N__11913\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__11913\,
            I => \Lab_UT.scdp.g0_0_i_1_1\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__11910\,
            I => \Lab_UT.scctrl.g1_1_1_1_cascade_\
        );

    \I__1881\ : InMux
    port map (
            O => \N__11907\,
            I => \N__11904\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__11904\,
            I => \Lab_UT.scctrl.g2_0\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__11901\,
            I => \N__11898\
        );

    \I__1878\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11895\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__11895\,
            I => \Lab_UT.scctrl.g1_3\
        );

    \I__1876\ : InMux
    port map (
            O => \N__11892\,
            I => \N__11889\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__11889\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__11886\,
            I => \N__11883\
        );

    \I__1873\ : InMux
    port map (
            O => \N__11883\,
            I => \N__11880\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__11880\,
            I => \N__11877\
        );

    \I__1871\ : Span4Mux_h
    port map (
            O => \N__11877\,
            I => \N__11874\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__11874\,
            I => \Lab_UT.scdp.byteToEncrypt_4\
        );

    \I__1869\ : InMux
    port map (
            O => \N__11871\,
            I => \N__11862\
        );

    \I__1868\ : InMux
    port map (
            O => \N__11870\,
            I => \N__11862\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11862\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__11862\,
            I => \N__11859\
        );

    \I__1865\ : Span4Mux_h
    port map (
            O => \N__11859\,
            I => \N__11856\
        );

    \I__1864\ : Odrv4
    port map (
            O => \N__11856\,
            I => \Lab_UT.scdp.b2a0.N_258_i\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11853\,
            I => \N__11850\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__11850\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1\
        );

    \I__1861\ : InMux
    port map (
            O => \N__11847\,
            I => \N__11842\
        );

    \I__1860\ : InMux
    port map (
            O => \N__11846\,
            I => \N__11837\
        );

    \I__1859\ : InMux
    port map (
            O => \N__11845\,
            I => \N__11834\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__11842\,
            I => \N__11831\
        );

    \I__1857\ : InMux
    port map (
            O => \N__11841\,
            I => \N__11827\
        );

    \I__1856\ : InMux
    port map (
            O => \N__11840\,
            I => \N__11824\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__11837\,
            I => \N__11817\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__11834\,
            I => \N__11817\
        );

    \I__1853\ : Span4Mux_v
    port map (
            O => \N__11831\,
            I => \N__11817\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11830\,
            I => \N__11814\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__11827\,
            I => \Lab_UT.scdp.d2eData_3_1_1\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__11824\,
            I => \Lab_UT.scdp.d2eData_3_1_1\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__11817\,
            I => \Lab_UT.scdp.d2eData_3_1_1\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__11814\,
            I => \Lab_UT.scdp.d2eData_3_1_1\
        );

    \I__1847\ : InMux
    port map (
            O => \N__11805\,
            I => \N__11802\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__11802\,
            I => \Lab_UT.scdp.d2eData_3_0_a2_0_4\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__11799\,
            I => \Lab_UT.scdp.d2eData_3_0_a2_0_4_cascade_\
        );

    \I__1844\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11793\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__11793\,
            I => \N__11788\
        );

    \I__1842\ : InMux
    port map (
            O => \N__11792\,
            I => \N__11783\
        );

    \I__1841\ : InMux
    port map (
            O => \N__11791\,
            I => \N__11783\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__11788\,
            I => \Lab_UT.scdp.N_246_i\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__11783\,
            I => \Lab_UT.scdp.N_246_i\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__11778\,
            I => \Lab_UT.scdp.N_246_i_cascade_\
        );

    \I__1837\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11772\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__11772\,
            I => \Lab_UT.scdp.u0.L4_tx_data_0_a2_1_6\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11766\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__11766\,
            I => \Lab_UT.scdp.N_256_i\
        );

    \I__1833\ : InMux
    port map (
            O => \N__11763\,
            I => \N__11759\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__11762\,
            I => \N__11756\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__11759\,
            I => \N__11753\
        );

    \I__1830\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11750\
        );

    \I__1829\ : Odrv12
    port map (
            O => \N__11753\,
            I => \Lab_UT.scdp.key0_2\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__11750\,
            I => \Lab_UT.scdp.key0_2\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__11745\,
            I => \Lab_UT.scdp.u1.g0_0_i_a5_0_0_1_cascade_\
        );

    \I__1826\ : InMux
    port map (
            O => \N__11742\,
            I => \N__11739\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__11739\,
            I => \Lab_UT.scdp.u1.g0_0_i_a5_0_2_1\
        );

    \I__1824\ : InMux
    port map (
            O => \N__11736\,
            I => \N__11733\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__11733\,
            I => \Lab_UT.scdp.N_6_1\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__11730\,
            I => \Lab_UT.scdp.d2eData_3_0_3_cascade_\
        );

    \I__1821\ : InMux
    port map (
            O => \N__11727\,
            I => \N__11721\
        );

    \I__1820\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11721\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__11721\,
            I => \Lab_UT.scdp.prng_lfsr_3\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__11718\,
            I => \N__11715\
        );

    \I__1817\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11712\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11712\,
            I => \N__11709\
        );

    \I__1815\ : Span4Mux_v
    port map (
            O => \N__11709\,
            I => \N__11706\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__11706\,
            I => \Lab_UT.scdp.byteToEncrypt_3\
        );

    \I__1813\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11700\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__11700\,
            I => \Lab_UT.scdp.d2eData_3_0_3\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__11697\,
            I => \N__11694\
        );

    \I__1810\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11687\
        );

    \I__1809\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11678\
        );

    \I__1808\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11678\
        );

    \I__1807\ : InMux
    port map (
            O => \N__11691\,
            I => \N__11678\
        );

    \I__1806\ : InMux
    port map (
            O => \N__11690\,
            I => \N__11678\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__11687\,
            I => \N__11673\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__11678\,
            I => \N__11673\
        );

    \I__1803\ : Span4Mux_v
    port map (
            O => \N__11673\,
            I => \N__11670\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__11670\,
            I => \Lab_UT.scdp.N_226_i\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11667\,
            I => \N__11664\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__11664\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__11661\,
            I => \N__11657\
        );

    \I__1798\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11652\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11648\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11643\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11655\,
            I => \N__11643\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__11652\,
            I => \N__11640\
        );

    \I__1793\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11637\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__11648\,
            I => \Lab_UT.scdp.d2eData_3_0_1\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__11643\,
            I => \Lab_UT.scdp.d2eData_3_0_1\
        );

    \I__1790\ : Odrv12
    port map (
            O => \N__11640\,
            I => \Lab_UT.scdp.d2eData_3_0_1\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__11637\,
            I => \Lab_UT.scdp.d2eData_3_0_1\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__11628\,
            I => \N__11624\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__11627\,
            I => \N__11618\
        );

    \I__1786\ : InMux
    port map (
            O => \N__11624\,
            I => \N__11612\
        );

    \I__1785\ : InMux
    port map (
            O => \N__11623\,
            I => \N__11612\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11607\
        );

    \I__1783\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11607\
        );

    \I__1782\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11604\
        );

    \I__1781\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11601\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11612\,
            I => \N__11598\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__11607\,
            I => \N__11593\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__11604\,
            I => \N__11593\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__11601\,
            I => \Lab_UT.scdp.u1.byteToDecrypt_1\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__11598\,
            I => \Lab_UT.scdp.u1.byteToDecrypt_1\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__11593\,
            I => \Lab_UT.scdp.u1.byteToDecrypt_1\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__11586\,
            I => \Lab_UT.scdp.u1.N_539_cascade_\
        );

    \I__1773\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11580\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__11580\,
            I => \N__11576\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11579\,
            I => \N__11571\
        );

    \I__1770\ : Span4Mux_v
    port map (
            O => \N__11576\,
            I => \N__11568\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11565\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11574\,
            I => \N__11562\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__11571\,
            I => \Lab_UT.scdp.N_255_i\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__11568\,
            I => \Lab_UT.scdp.N_255_i\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__11565\,
            I => \Lab_UT.scdp.N_255_i\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__11562\,
            I => \Lab_UT.scdp.N_255_i\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11553\,
            I => \N__11549\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11552\,
            I => \N__11541\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__11549\,
            I => \N__11538\
        );

    \I__1760\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11529\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11529\
        );

    \I__1758\ : InMux
    port map (
            O => \N__11546\,
            I => \N__11529\
        );

    \I__1757\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11529\
        );

    \I__1756\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11526\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__11541\,
            I => \Lab_UT.scdp.N_228_i\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__11538\,
            I => \Lab_UT.scdp.N_228_i\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__11529\,
            I => \Lab_UT.scdp.N_228_i\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__11526\,
            I => \Lab_UT.scdp.N_228_i\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__11517\,
            I => \Lab_UT.scdp.N_426_cascade_\
        );

    \I__1750\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11511\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__11511\,
            I => \N__11508\
        );

    \I__1748\ : Sp12to4
    port map (
            O => \N__11508\,
            I => \N__11505\
        );

    \I__1747\ : Odrv12
    port map (
            O => \N__11505\,
            I => \Lab_UT.scdp.q_RNI47LGA_1\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11499\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__11499\,
            I => \Lab_UT.scdp.N_73\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__11496\,
            I => \Lab_UT.scdp.N_73_cascade_\
        );

    \I__1743\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11490\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__11490\,
            I => \N__11487\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__11487\,
            I => \Lab_UT.scctrl.delayload\
        );

    \I__1740\ : InMux
    port map (
            O => \N__11484\,
            I => \N__11481\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__11481\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__11478\,
            I => \N__11475\
        );

    \I__1737\ : InMux
    port map (
            O => \N__11475\,
            I => \N__11472\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11472\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11466\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__11466\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__11463\,
            I => \Lab_UT.scdp.d2eData_3_5_cascade_\
        );

    \I__1732\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11456\
        );

    \I__1731\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11453\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__11456\,
            I => \N__11450\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__11453\,
            I => \Lab_UT.scdp.N_225_i_1\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__11450\,
            I => \Lab_UT.scdp.N_225_i_1\
        );

    \I__1727\ : InMux
    port map (
            O => \N__11445\,
            I => \N__11442\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__11442\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__11439\,
            I => \buart.Z_rx.N_230_cascade_\
        );

    \I__1724\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11433\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__11433\,
            I => \N__11429\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__11432\,
            I => \N__11426\
        );

    \I__1721\ : Span4Mux_h
    port map (
            O => \N__11429\,
            I => \N__11423\
        );

    \I__1720\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11420\
        );

    \I__1719\ : Odrv4
    port map (
            O => \N__11423\,
            I => \Lab_UT.scdp.key0_7\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__11420\,
            I => \Lab_UT.scdp.key0_7\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11415\,
            I => \N__11412\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__11412\,
            I => \N__11409\
        );

    \I__1715\ : Span4Mux_v
    port map (
            O => \N__11409\,
            I => \N__11405\
        );

    \I__1714\ : InMux
    port map (
            O => \N__11408\,
            I => \N__11402\
        );

    \I__1713\ : Odrv4
    port map (
            O => \N__11405\,
            I => \Lab_UT.scdp.key0_3\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__11402\,
            I => \Lab_UT.scdp.key0_3\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__11397\,
            I => \Lab_UT.scdp.binVal_2_cascade_\
        );

    \I__1710\ : CascadeMux
    port map (
            O => \N__11394\,
            I => \Lab_UT.scctrl.g1_0_1_cascade_\
        );

    \I__1709\ : InMux
    port map (
            O => \N__11391\,
            I => \N__11388\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__11388\,
            I => \N__11385\
        );

    \I__1707\ : Span4Mux_v
    port map (
            O => \N__11385\,
            I => \N__11381\
        );

    \I__1706\ : InMux
    port map (
            O => \N__11384\,
            I => \N__11378\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__11381\,
            I => \Lab_UT.scdp.N_276\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__11378\,
            I => \Lab_UT.scdp.N_276\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__11373\,
            I => \N__11370\
        );

    \I__1702\ : InMux
    port map (
            O => \N__11370\,
            I => \N__11367\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__11367\,
            I => \N__11364\
        );

    \I__1700\ : Span4Mux_h
    port map (
            O => \N__11364\,
            I => \N__11361\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__11361\,
            I => \Lab_UT.scdp.msBitsi.N_41\
        );

    \I__1698\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11355\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__11355\,
            I => \N__11352\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__11352\,
            I => \N__11349\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__11349\,
            I => \ufifo.txdataDZ0Z_0\
        );

    \I__1694\ : InMux
    port map (
            O => \N__11346\,
            I => \N__11343\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__11343\,
            I => \Lab_UT.scctrl.N_46\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__11340\,
            I => \N__11337\
        );

    \I__1691\ : InMux
    port map (
            O => \N__11337\,
            I => \N__11334\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__11334\,
            I => \N__11331\
        );

    \I__1689\ : Span4Mux_s2_h
    port map (
            O => \N__11331\,
            I => \N__11328\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__11328\,
            I => \buart.Z_rx.sample_i_0_a2_0\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__11325\,
            I => \N__11321\
        );

    \I__1686\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11318\
        );

    \I__1685\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11315\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__11318\,
            I => \N__11312\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__11315\,
            I => \buart.Z_rx.N_230\
        );

    \I__1682\ : Odrv12
    port map (
            O => \N__11312\,
            I => \buart.Z_rx.N_230\
        );

    \I__1681\ : SRMux
    port map (
            O => \N__11307\,
            I => \N__11304\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__11304\,
            I => \N__11298\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__11303\,
            I => \N__11295\
        );

    \I__1678\ : CEMux
    port map (
            O => \N__11302\,
            I => \N__11292\
        );

    \I__1677\ : InMux
    port map (
            O => \N__11301\,
            I => \N__11289\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__11298\,
            I => \N__11286\
        );

    \I__1675\ : InMux
    port map (
            O => \N__11295\,
            I => \N__11283\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__11292\,
            I => \N__11280\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__11289\,
            I => \N__11277\
        );

    \I__1672\ : IoSpan4Mux
    port map (
            O => \N__11286\,
            I => \N__11272\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__11283\,
            I => \N__11272\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__11280\,
            I => \N__11269\
        );

    \I__1669\ : Span4Mux_s1_h
    port map (
            O => \N__11277\,
            I => \N__11264\
        );

    \I__1668\ : Span4Mux_s1_h
    port map (
            O => \N__11272\,
            I => \N__11264\
        );

    \I__1667\ : Span4Mux_s2_h
    port map (
            O => \N__11269\,
            I => \N__11261\
        );

    \I__1666\ : Span4Mux_h
    port map (
            O => \N__11264\,
            I => \N__11258\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__11261\,
            I => \ufifo.txDataValidDZ0\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__11258\,
            I => \ufifo.txDataValidDZ0\
        );

    \I__1663\ : InMux
    port map (
            O => \N__11253\,
            I => \N__11250\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__11250\,
            I => \N__11246\
        );

    \I__1661\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11243\
        );

    \I__1660\ : Span4Mux_v
    port map (
            O => \N__11246\,
            I => \N__11238\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__11243\,
            I => \N__11238\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__11238\,
            I => \N_233_reti\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__11235\,
            I => \Lab_UT.scctrl.g1_0_1_0_cascade_\
        );

    \I__1656\ : InMux
    port map (
            O => \N__11232\,
            I => \N__11225\
        );

    \I__1655\ : InMux
    port map (
            O => \N__11231\,
            I => \N__11225\
        );

    \I__1654\ : InMux
    port map (
            O => \N__11230\,
            I => \N__11222\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__11225\,
            I => \Lab_UT.sccElsBitsLd\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__11222\,
            I => \Lab_UT.sccElsBitsLd\
        );

    \I__1651\ : CEMux
    port map (
            O => \N__11217\,
            I => \N__11213\
        );

    \I__1650\ : CEMux
    port map (
            O => \N__11216\,
            I => \N__11210\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__11213\,
            I => \N__11207\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__11210\,
            I => \N__11204\
        );

    \I__1647\ : Span4Mux_v
    port map (
            O => \N__11207\,
            I => \N__11201\
        );

    \I__1646\ : Span4Mux_h
    port map (
            O => \N__11204\,
            I => \N__11198\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__11201\,
            I => \Lab_UT.scdp.sccElsBitsLd_0\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__11198\,
            I => \Lab_UT.scdp.sccElsBitsLd_0\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11190\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__11190\,
            I => \N__11187\
        );

    \I__1641\ : Span4Mux_h
    port map (
            O => \N__11187\,
            I => \N__11184\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__11184\,
            I => \Lab_UT.scdp.msBitsi.q_esr_RNI679EZ0Z_6\
        );

    \I__1639\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11178\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__11178\,
            I => \N__11175\
        );

    \I__1637\ : Odrv12
    port map (
            O => \N__11175\,
            I => \ufifo.txdataDZ0Z_6\
        );

    \I__1636\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11169\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__11169\,
            I => \Lab_UT.scctrl.N_534\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__11166\,
            I => \Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0_cascade_\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11160\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__11160\,
            I => \Lab_UT.scctrl.N_415_0\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__11157\,
            I => \N__11154\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11154\,
            I => \N__11151\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__11151\,
            I => \Lab_UT.scctrl.g1_0_0\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__11148\,
            I => \Lab_UT.scctrl.g1_0_2_cascade_\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__11145\,
            I => \Lab_UT.scctrl.next_state_0_0_2_cascade_\
        );

    \I__1626\ : InMux
    port map (
            O => \N__11142\,
            I => \N__11139\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__11139\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11136\,
            I => \N__11133\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__11133\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30\
        );

    \I__1622\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11127\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__11127\,
            I => \N__11124\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__11124\,
            I => \resetGen.N_243\
        );

    \I__1619\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11118\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__11118\,
            I => \N__11115\
        );

    \I__1617\ : Span4Mux_v
    port map (
            O => \N__11115\,
            I => \N__11112\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__11112\,
            I => \buart.bu_rx_data_i_2_4\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__11109\,
            I => \N__11105\
        );

    \I__1614\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11100\
        );

    \I__1613\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11100\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__11100\,
            I => \Lab_UT.scdp.N_225_i_0\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__11097\,
            I => \Lab_UT.scdp.u1.g0_0_i_a5_0_2_cascade_\
        );

    \I__1610\ : InMux
    port map (
            O => \N__11094\,
            I => \N__11091\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__11091\,
            I => \Lab_UT.scdp.N_6\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__11088\,
            I => \Lab_UT.scdp.u1.g0_0_i_a5_0_2_0_cascade_\
        );

    \I__1607\ : InMux
    port map (
            O => \N__11085\,
            I => \N__11082\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__11082\,
            I => \Lab_UT.scdp.N_6_0\
        );

    \I__1605\ : InMux
    port map (
            O => \N__11079\,
            I => \N__11076\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__11076\,
            I => \N__11071\
        );

    \I__1603\ : InMux
    port map (
            O => \N__11075\,
            I => \N__11066\
        );

    \I__1602\ : InMux
    port map (
            O => \N__11074\,
            I => \N__11066\
        );

    \I__1601\ : Odrv12
    port map (
            O => \N__11071\,
            I => \Lab_UT.scdp.d2eData_3_0_a2_0_6\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__11066\,
            I => \Lab_UT.scdp.d2eData_3_0_a2_0_6\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__11061\,
            I => \N__11056\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__11060\,
            I => \N__11053\
        );

    \I__1597\ : InMux
    port map (
            O => \N__11059\,
            I => \N__11050\
        );

    \I__1596\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11045\
        );

    \I__1595\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11045\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__11050\,
            I => \N__11042\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__11045\,
            I => \N__11039\
        );

    \I__1592\ : Odrv12
    port map (
            O => \N__11042\,
            I => \Lab_UT.scdp.prng_lfsr_14\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__11039\,
            I => \Lab_UT.scdp.prng_lfsr_14\
        );

    \I__1590\ : InMux
    port map (
            O => \N__11034\,
            I => \N__11031\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__11031\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17\
        );

    \I__1588\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11025\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__11025\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__11022\,
            I => \N__11019\
        );

    \I__1585\ : InMux
    port map (
            O => \N__11019\,
            I => \N__11016\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__11016\,
            I => \N__11013\
        );

    \I__1583\ : Odrv4
    port map (
            O => \N__11013\,
            I => \Lab_UT.scdp.msBitsi.N_1919_0\
        );

    \I__1582\ : InMux
    port map (
            O => \N__11010\,
            I => \N__11007\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__11007\,
            I => \N__11004\
        );

    \I__1580\ : Sp12to4
    port map (
            O => \N__11004\,
            I => \N__11001\
        );

    \I__1579\ : Odrv12
    port map (
            O => \N__11001\,
            I => \ufifo.txdataDZ0Z_2\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__10998\,
            I => \N__10995\
        );

    \I__1577\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10992\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__10992\,
            I => \N__10989\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__10989\,
            I => \Lab_UT.scdp.msBitsi.N_1917_0\
        );

    \I__1574\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10983\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__10983\,
            I => \N__10980\
        );

    \I__1572\ : Span4Mux_v
    port map (
            O => \N__10980\,
            I => \N__10977\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__10977\,
            I => \ufifo.txdataDZ0Z_4\
        );

    \I__1570\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10971\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__10971\,
            I => \Lab_UT.scdp.N_552\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__10968\,
            I => \Lab_UT.scdp.N_228_i_0_cascade_\
        );

    \I__1567\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10959\
        );

    \I__1566\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10959\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__10959\,
            I => \N__10956\
        );

    \I__1564\ : Odrv12
    port map (
            O => \N__10956\,
            I => \Lab_UT.scdp.u0.byteToDecrypt_6\
        );

    \I__1563\ : InMux
    port map (
            O => \N__10953\,
            I => \N__10950\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__10950\,
            I => \N__10947\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__10947\,
            I => \N__10944\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__10944\,
            I => \Lab_UT.scdp.lfsrInst.N_234_i_0\
        );

    \I__1559\ : InMux
    port map (
            O => \N__10941\,
            I => \N__10938\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__10938\,
            I => \Lab_UT.scdp.g0_0_i_1\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__10935\,
            I => \Lab_UT.scdp.d2eData_3_0_1_cascade_\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10932\,
            I => \N__10929\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__10929\,
            I => \Lab_UT.scdp.msBitsi.msBitsD_1\
        );

    \I__1554\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10923\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__10923\,
            I => \N__10920\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__10920\,
            I => \Lab_UT.scdp.lsBitsD_1\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__10917\,
            I => \Lab_UT.scdp.msBitsi.N_43_cascade_\
        );

    \I__1550\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10911\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__10911\,
            I => \N__10908\
        );

    \I__1548\ : Span4Mux_v
    port map (
            O => \N__10908\,
            I => \N__10905\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__10905\,
            I => \ufifo.txdataDZ0Z_1\
        );

    \I__1546\ : InMux
    port map (
            O => \N__10902\,
            I => \N__10899\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__10899\,
            I => \Lab_UT.scdp.msBitsi.msBitsD_2\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10893\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__10893\,
            I => \N__10890\
        );

    \I__1542\ : Span4Mux_v
    port map (
            O => \N__10890\,
            I => \N__10887\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__10887\,
            I => \Lab_UT.scdp.lsBitsD_2\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10881\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__10881\,
            I => \Lab_UT.scdp.msBitsi.msBitsD_4\
        );

    \I__1538\ : InMux
    port map (
            O => \N__10878\,
            I => \N__10875\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__10875\,
            I => \N__10872\
        );

    \I__1536\ : Odrv12
    port map (
            O => \N__10872\,
            I => \Lab_UT.scdp.lsBitsD_4\
        );

    \I__1535\ : InMux
    port map (
            O => \N__10869\,
            I => \N__10866\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__10866\,
            I => \N__10863\
        );

    \I__1533\ : Span4Mux_v
    port map (
            O => \N__10863\,
            I => \N__10859\
        );

    \I__1532\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10856\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__10859\,
            I => \Lab_UT.scdp.lsBitsi.lsBitsDZ0Z_5\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__10856\,
            I => \Lab_UT.scdp.lsBitsi.lsBitsDZ0Z_5\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__10851\,
            I => \Lab_UT.scdp.N_332_i_1_cascade_\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10845\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__10845\,
            I => \N__10842\
        );

    \I__1526\ : Span4Mux_v
    port map (
            O => \N__10842\,
            I => \N__10839\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__10839\,
            I => \ufifo.txdataDZ0Z_5\
        );

    \I__1524\ : InMux
    port map (
            O => \N__10836\,
            I => \N__10833\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__10833\,
            I => \N__10824\
        );

    \I__1522\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10813\
        );

    \I__1521\ : InMux
    port map (
            O => \N__10831\,
            I => \N__10813\
        );

    \I__1520\ : InMux
    port map (
            O => \N__10830\,
            I => \N__10813\
        );

    \I__1519\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10813\
        );

    \I__1518\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10813\
        );

    \I__1517\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10810\
        );

    \I__1516\ : Span4Mux_h
    port map (
            O => \N__10824\,
            I => \N__10807\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__10813\,
            I => \N__10804\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__10810\,
            I => \Lab_UT.sccEmsBitsSl\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__10807\,
            I => \Lab_UT.sccEmsBitsSl\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__10804\,
            I => \Lab_UT.sccEmsBitsSl\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__10797\,
            I => \N__10794\
        );

    \I__1510\ : InMux
    port map (
            O => \N__10794\,
            I => \N__10791\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10791\,
            I => \Lab_UT.scdp.msBitsi.msBitsD_3\
        );

    \I__1508\ : InMux
    port map (
            O => \N__10788\,
            I => \N__10784\
        );

    \I__1507\ : InMux
    port map (
            O => \N__10787\,
            I => \N__10781\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__10784\,
            I => \N__10778\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__10781\,
            I => \Lab_UT.scdp.lsBitsD_3\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__10778\,
            I => \Lab_UT.scdp.lsBitsD_3\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10770\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__10770\,
            I => \N__10767\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__10767\,
            I => \Lab_UT.scdp.g0_0_i_1_0\
        );

    \I__1500\ : InMux
    port map (
            O => \N__10764\,
            I => \N__10761\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__10761\,
            I => \Lab_UT.scdp.msBitsi.N_1915_0\
        );

    \I__1498\ : InMux
    port map (
            O => \N__10758\,
            I => \N__10755\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__10755\,
            I => \N__10752\
        );

    \I__1496\ : Span4Mux_h
    port map (
            O => \N__10752\,
            I => \N__10749\
        );

    \I__1495\ : Span4Mux_v
    port map (
            O => \N__10749\,
            I => \N__10746\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__10746\,
            I => \ufifo.txdataDZ0Z_3\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__10743\,
            I => \N__10740\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10737\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__10737\,
            I => \N__10734\
        );

    \I__1490\ : Span4Mux_h
    port map (
            O => \N__10734\,
            I => \N__10731\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__10731\,
            I => \Lab_UT.scdp.byteToEncrypt_6\
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__10728\,
            I => \Lab_UT.scdp.b2a0.N_238_i_cascade_\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__10725\,
            I => \N__10719\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__10724\,
            I => \N__10716\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10704\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10722\,
            I => \N__10704\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10719\,
            I => \N__10704\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10716\,
            I => \N__10704\
        );

    \I__1481\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10704\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__10704\,
            I => \Lab_UT.scdp.b2a0.N_238_i\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__10701\,
            I => \N__10697\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__10700\,
            I => \N__10690\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10685\
        );

    \I__1476\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10685\
        );

    \I__1475\ : InMux
    port map (
            O => \N__10695\,
            I => \N__10676\
        );

    \I__1474\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10676\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10693\,
            I => \N__10676\
        );

    \I__1472\ : InMux
    port map (
            O => \N__10690\,
            I => \N__10676\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__10685\,
            I => \N__10671\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__10676\,
            I => \N__10671\
        );

    \I__1469\ : Span4Mux_h
    port map (
            O => \N__10671\,
            I => \N__10668\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__10668\,
            I => \Lab_UT.scdp.b2a0.N_227_i\
        );

    \I__1467\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10662\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__10662\,
            I => \N__10659\
        );

    \I__1465\ : Span4Mux_h
    port map (
            O => \N__10659\,
            I => \N__10656\
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__10656\,
            I => \Lab_UT.scdp.msBitsi.msBitsD_6\
        );

    \I__1463\ : InMux
    port map (
            O => \N__10653\,
            I => \N__10646\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10646\
        );

    \I__1461\ : InMux
    port map (
            O => \N__10651\,
            I => \N__10643\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10638\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__10643\,
            I => \N__10638\
        );

    \I__1458\ : Span4Mux_h
    port map (
            O => \N__10638\,
            I => \N__10635\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__10635\,
            I => \Lab_UT.scdp.byteToEncrypt_5\
        );

    \I__1456\ : InMux
    port map (
            O => \N__10632\,
            I => \N__10620\
        );

    \I__1455\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10620\
        );

    \I__1454\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10620\
        );

    \I__1453\ : InMux
    port map (
            O => \N__10629\,
            I => \N__10620\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__10620\,
            I => \Lab_UT.scdp.b2a0.N_224_i\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10617\,
            I => \N__10614\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__10614\,
            I => \Lab_UT.scdp.msBitsi.msBitsD_0\
        );

    \I__1449\ : InMux
    port map (
            O => \N__10611\,
            I => \N__10608\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__10608\,
            I => \N__10605\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__10605\,
            I => \Lab_UT.scdp.lsBitsD_0\
        );

    \I__1446\ : InMux
    port map (
            O => \N__10602\,
            I => \N__10599\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__10599\,
            I => \N__10596\
        );

    \I__1444\ : Span4Mux_h
    port map (
            O => \N__10596\,
            I => \N__10593\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__10593\,
            I => \Lab_UT.scdp.byteToEncrypt_1\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__10590\,
            I => \N__10585\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__10589\,
            I => \N__10581\
        );

    \I__1440\ : InMux
    port map (
            O => \N__10588\,
            I => \N__10572\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10585\,
            I => \N__10572\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10584\,
            I => \N__10572\
        );

    \I__1437\ : InMux
    port map (
            O => \N__10581\,
            I => \N__10572\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__10572\,
            I => \N__10569\
        );

    \I__1435\ : Span4Mux_h
    port map (
            O => \N__10569\,
            I => \N__10566\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__10566\,
            I => \Lab_UT.scdp.byteToEncrypt_2\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__10563\,
            I => \Lab_UT.scdp.b2a1.N_220_i_cascade_\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__10560\,
            I => \N__10557\
        );

    \I__1431\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10545\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10545\
        );

    \I__1429\ : InMux
    port map (
            O => \N__10555\,
            I => \N__10545\
        );

    \I__1428\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10545\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__10545\,
            I => \Lab_UT.scdp.b2a1.N_220_i\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__10542\,
            I => \Lab_UT.scdp.N_282_cascade_\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10533\
        );

    \I__1424\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10533\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__10533\,
            I => \Lab_UT.scdp.b2a1.N_293\
        );

    \I__1422\ : IoInMux
    port map (
            O => \N__10530\,
            I => \N__10527\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__10527\,
            I => \N__10523\
        );

    \I__1420\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10520\
        );

    \I__1419\ : Span4Mux_s3_v
    port map (
            O => \N__10523\,
            I => \N__10517\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__10520\,
            I => \N__10512\
        );

    \I__1417\ : Span4Mux_v
    port map (
            O => \N__10517\,
            I => \N__10512\
        );

    \I__1416\ : Odrv4
    port map (
            O => \N__10512\,
            I => \Lab_UT.scctrl.sccLdLFSR\
        );

    \I__1415\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10506\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__10506\,
            I => \Lab_UT.scctrl.EmsLoaded\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__10503\,
            I => \Lab_UT.scctrl.EmsLoaded_cascade_\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__10500\,
            I => \Lab_UT.sccElsBitsLd_cascade_\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10497\,
            I => \N__10494\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__10494\,
            I => \Lab_UT.scdp.lsBits_i_1_6\
        );

    \I__1409\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10487\
        );

    \I__1408\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10484\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__10487\,
            I => \N__10481\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__10484\,
            I => \Lab_UT.scdp.lsBitsD_6\
        );

    \I__1405\ : Odrv4
    port map (
            O => \N__10481\,
            I => \Lab_UT.scdp.lsBitsD_6\
        );

    \I__1404\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10472\
        );

    \I__1403\ : InMux
    port map (
            O => \N__10475\,
            I => \N__10469\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__10472\,
            I => \Lab_UT.scdp.N_282\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__10469\,
            I => \Lab_UT.scdp.N_282\
        );

    \I__1400\ : InMux
    port map (
            O => \N__10464\,
            I => \N__10458\
        );

    \I__1399\ : InMux
    port map (
            O => \N__10463\,
            I => \N__10458\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__10458\,
            I => \N__10455\
        );

    \I__1397\ : Odrv12
    port map (
            O => \N__10455\,
            I => \resetGen.N_274\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10446\
        );

    \I__1395\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10446\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__10446\,
            I => \N__10441\
        );

    \I__1393\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10436\
        );

    \I__1392\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10436\
        );

    \I__1391\ : Odrv12
    port map (
            O => \N__10441\,
            I => \resetGen.N_421\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__10436\,
            I => \resetGen.N_421\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__10431\,
            I => \N__10427\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__10430\,
            I => \N__10424\
        );

    \I__1387\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10419\
        );

    \I__1386\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10419\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__10419\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__1384\ : InMux
    port map (
            O => \N__10416\,
            I => \N__10413\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__10413\,
            I => \N__10409\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__10412\,
            I => \N__10406\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__10409\,
            I => \N__10397\
        );

    \I__1380\ : InMux
    port map (
            O => \N__10406\,
            I => \N__10394\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10389\
        );

    \I__1378\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10389\
        );

    \I__1377\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10384\
        );

    \I__1376\ : InMux
    port map (
            O => \N__10402\,
            I => \N__10384\
        );

    \I__1375\ : InMux
    port map (
            O => \N__10401\,
            I => \N__10381\
        );

    \I__1374\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10378\
        );

    \I__1373\ : Sp12to4
    port map (
            O => \N__10397\,
            I => \N__10375\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__10394\,
            I => \N__10372\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__10389\,
            I => \N__10369\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__10384\,
            I => ufifo_tx_fsm_cstate_0
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__10381\,
            I => ufifo_tx_fsm_cstate_0
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__10378\,
            I => ufifo_tx_fsm_cstate_0
        );

    \I__1367\ : Odrv12
    port map (
            O => \N__10375\,
            I => ufifo_tx_fsm_cstate_0
        );

    \I__1366\ : Odrv4
    port map (
            O => \N__10372\,
            I => ufifo_tx_fsm_cstate_0
        );

    \I__1365\ : Odrv12
    port map (
            O => \N__10369\,
            I => ufifo_tx_fsm_cstate_0
        );

    \I__1364\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10353\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__10353\,
            I => \N__10350\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__10350\,
            I => \ufifo.fifo.fifo_txdata_0\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__10347\,
            I => \N__10344\
        );

    \I__1360\ : InMux
    port map (
            O => \N__10344\,
            I => \N__10338\
        );

    \I__1359\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10338\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__10338\,
            I => \N__10335\
        );

    \I__1357\ : Span4Mux_h
    port map (
            O => \N__10335\,
            I => \N__10332\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__10332\,
            I => \Lab_UT.scdp.byteToEncrypt_0\
        );

    \I__1355\ : InMux
    port map (
            O => \N__10329\,
            I => \ufifo.fifo.un1_rdaddr_cry_5\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__10326\,
            I => \N__10323\
        );

    \I__1353\ : InMux
    port map (
            O => \N__10323\,
            I => \N__10318\
        );

    \I__1352\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10315\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10312\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__10318\,
            I => \N__10307\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__10315\,
            I => \N__10307\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__10312\,
            I => \N__10302\
        );

    \I__1347\ : Span4Mux_v
    port map (
            O => \N__10307\,
            I => \N__10302\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__10302\,
            I => \ufifo.fifo.rdaddrZ0Z_7\
        );

    \I__1345\ : InMux
    port map (
            O => \N__10299\,
            I => \ufifo.fifo.un1_rdaddr_cry_6\
        );

    \I__1344\ : InMux
    port map (
            O => \N__10296\,
            I => \bfn_4_5_0_\
        );

    \I__1343\ : CascadeMux
    port map (
            O => \N__10293\,
            I => \N__10289\
        );

    \I__1342\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10285\
        );

    \I__1341\ : InMux
    port map (
            O => \N__10289\,
            I => \N__10282\
        );

    \I__1340\ : InMux
    port map (
            O => \N__10288\,
            I => \N__10279\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__10285\,
            I => \N__10276\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__10282\,
            I => \ufifo.fifo.rdaddrZ0Z_8\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__10279\,
            I => \ufifo.fifo.rdaddrZ0Z_8\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__10276\,
            I => \ufifo.fifo.rdaddrZ0Z_8\
        );

    \I__1335\ : InMux
    port map (
            O => \N__10269\,
            I => \N__10264\
        );

    \I__1334\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10259\
        );

    \I__1333\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10259\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10256\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__10259\,
            I => \N__10253\
        );

    \I__1330\ : Span4Mux_s3_h
    port map (
            O => \N__10256\,
            I => \N__10250\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__10253\,
            I => \N_251\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__10250\,
            I => \N_251\
        );

    \I__1327\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10242\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__10242\,
            I => \ufifo.fifo.fifo_txdata_1\
        );

    \I__1325\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10236\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__10236\,
            I => \N__10233\
        );

    \I__1323\ : Span4Mux_v
    port map (
            O => \N__10233\,
            I => \N__10230\
        );

    \I__1322\ : Odrv4
    port map (
            O => \N__10230\,
            I => \ufifo.sb_ram512x8_inst_RNIKRN11\
        );

    \I__1321\ : InMux
    port map (
            O => \N__10227\,
            I => \N__10224\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__10224\,
            I => \N__10220\
        );

    \I__1319\ : InMux
    port map (
            O => \N__10223\,
            I => \N__10217\
        );

    \I__1318\ : Span4Mux_s3_h
    port map (
            O => \N__10220\,
            I => \N__10214\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__10217\,
            I => \N__10211\
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__10214\,
            I => ufifo_fifo_txdata_rdy
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__10211\,
            I => ufifo_fifo_txdata_rdy
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__10206\,
            I => \N__10202\
        );

    \I__1313\ : InMux
    port map (
            O => \N__10205\,
            I => \N__10199\
        );

    \I__1312\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10196\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__10199\,
            I => \N__10193\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__10196\,
            I => \N__10190\
        );

    \I__1309\ : Span4Mux_s3_h
    port map (
            O => \N__10193\,
            I => \N__10187\
        );

    \I__1308\ : Odrv12
    port map (
            O => \N__10190\,
            I => \buart.Z_tx.N_278\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__10187\,
            I => \buart.Z_tx.N_278\
        );

    \I__1306\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10170\
        );

    \I__1305\ : InMux
    port map (
            O => \N__10181\,
            I => \N__10170\
        );

    \I__1304\ : InMux
    port map (
            O => \N__10180\,
            I => \N__10170\
        );

    \I__1303\ : InMux
    port map (
            O => \N__10179\,
            I => \N__10170\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__10170\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__10167\,
            I => \N__10164\
        );

    \I__1300\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10155\
        );

    \I__1299\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10155\
        );

    \I__1298\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10155\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__10155\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__1296\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10148\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10151\,
            I => \N__10145\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__10148\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__10145\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1292\ : CEMux
    port map (
            O => \N__10140\,
            I => \N__10136\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__10139\,
            I => \N__10131\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__10136\,
            I => \N__10127\
        );

    \I__1289\ : InMux
    port map (
            O => \N__10135\,
            I => \N__10124\
        );

    \I__1288\ : InMux
    port map (
            O => \N__10134\,
            I => \N__10121\
        );

    \I__1287\ : InMux
    port map (
            O => \N__10131\,
            I => \N__10118\
        );

    \I__1286\ : SRMux
    port map (
            O => \N__10130\,
            I => \N__10115\
        );

    \I__1285\ : Span4Mux_v
    port map (
            O => \N__10127\,
            I => \N__10112\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10109\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__10121\,
            I => \N__10104\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__10118\,
            I => \N__10104\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__10115\,
            I => \N__10099\
        );

    \I__1280\ : Span4Mux_s2_h
    port map (
            O => \N__10112\,
            I => \N__10099\
        );

    \I__1279\ : Span4Mux_h
    port map (
            O => \N__10109\,
            I => \N__10096\
        );

    \I__1278\ : Span4Mux_h
    port map (
            O => \N__10104\,
            I => \N__10093\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__10099\,
            I => \ufifo.popFifo\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__10096\,
            I => \ufifo.popFifo\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__10093\,
            I => \ufifo.popFifo\
        );

    \I__1274\ : CascadeMux
    port map (
            O => \N__10086\,
            I => \N__10082\
        );

    \I__1273\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10079\
        );

    \I__1272\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10076\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__10079\,
            I => \N__10072\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__10076\,
            I => \N__10069\
        );

    \I__1269\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10066\
        );

    \I__1268\ : Span4Mux_s3_h
    port map (
            O => \N__10072\,
            I => \N__10063\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__10069\,
            I => \ufifo.fifo.rdaddrZ0Z_0\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__10066\,
            I => \ufifo.fifo.rdaddrZ0Z_0\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__10063\,
            I => \ufifo.fifo.rdaddrZ0Z_0\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__10056\,
            I => \N__10053\
        );

    \I__1263\ : InMux
    port map (
            O => \N__10053\,
            I => \N__10050\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__10050\,
            I => \N__10046\
        );

    \I__1261\ : InMux
    port map (
            O => \N__10049\,
            I => \N__10043\
        );

    \I__1260\ : Span4Mux_v
    port map (
            O => \N__10046\,
            I => \N__10037\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__10043\,
            I => \N__10037\
        );

    \I__1258\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10034\
        );

    \I__1257\ : Span4Mux_s3_h
    port map (
            O => \N__10037\,
            I => \N__10031\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__10034\,
            I => \ufifo.fifo.rdaddrZ0Z_1\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__10031\,
            I => \ufifo.fifo.rdaddrZ0Z_1\
        );

    \I__1254\ : InMux
    port map (
            O => \N__10026\,
            I => \ufifo.fifo.un1_rdaddr_cry_0\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__10023\,
            I => \N__10019\
        );

    \I__1252\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10016\
        );

    \I__1251\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10013\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__10016\,
            I => \N__10009\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__10013\,
            I => \N__10006\
        );

    \I__1248\ : InMux
    port map (
            O => \N__10012\,
            I => \N__10003\
        );

    \I__1247\ : Span4Mux_s3_h
    port map (
            O => \N__10009\,
            I => \N__10000\
        );

    \I__1246\ : Odrv4
    port map (
            O => \N__10006\,
            I => \ufifo.fifo.rdaddrZ0Z_2\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__10003\,
            I => \ufifo.fifo.rdaddrZ0Z_2\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__10000\,
            I => \ufifo.fifo.rdaddrZ0Z_2\
        );

    \I__1243\ : InMux
    port map (
            O => \N__9993\,
            I => \ufifo.fifo.un1_rdaddr_cry_1\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__9990\,
            I => \N__9987\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9987\,
            I => \N__9983\
        );

    \I__1240\ : InMux
    port map (
            O => \N__9986\,
            I => \N__9980\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__9983\,
            I => \N__9976\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__9980\,
            I => \N__9973\
        );

    \I__1237\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9970\
        );

    \I__1236\ : Span4Mux_v
    port map (
            O => \N__9976\,
            I => \N__9965\
        );

    \I__1235\ : Span4Mux_s3_h
    port map (
            O => \N__9973\,
            I => \N__9965\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__9970\,
            I => \ufifo.fifo.rdaddrZ0Z_3\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__9965\,
            I => \ufifo.fifo.rdaddrZ0Z_3\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9960\,
            I => \ufifo.fifo.un1_rdaddr_cry_2\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__9957\,
            I => \N__9954\
        );

    \I__1230\ : InMux
    port map (
            O => \N__9954\,
            I => \N__9950\
        );

    \I__1229\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9947\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__9950\,
            I => \N__9941\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__9947\,
            I => \N__9941\
        );

    \I__1226\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9938\
        );

    \I__1225\ : Span4Mux_s3_h
    port map (
            O => \N__9941\,
            I => \N__9935\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__9938\,
            I => \ufifo.fifo.rdaddrZ0Z_4\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__9935\,
            I => \ufifo.fifo.rdaddrZ0Z_4\
        );

    \I__1222\ : InMux
    port map (
            O => \N__9930\,
            I => \ufifo.fifo.un1_rdaddr_cry_3\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__9927\,
            I => \N__9923\
        );

    \I__1220\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9920\
        );

    \I__1219\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9916\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__9920\,
            I => \N__9913\
        );

    \I__1217\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9910\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__9916\,
            I => \N__9905\
        );

    \I__1215\ : Span4Mux_s3_h
    port map (
            O => \N__9913\,
            I => \N__9905\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__9910\,
            I => \ufifo.fifo.rdaddrZ0Z_5\
        );

    \I__1213\ : Odrv4
    port map (
            O => \N__9905\,
            I => \ufifo.fifo.rdaddrZ0Z_5\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9900\,
            I => \ufifo.fifo.un1_rdaddr_cry_4\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__9897\,
            I => \N__9894\
        );

    \I__1210\ : InMux
    port map (
            O => \N__9894\,
            I => \N__9890\
        );

    \I__1209\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9887\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__9890\,
            I => \N__9883\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__9887\,
            I => \N__9880\
        );

    \I__1206\ : InMux
    port map (
            O => \N__9886\,
            I => \N__9877\
        );

    \I__1205\ : Span4Mux_s3_h
    port map (
            O => \N__9883\,
            I => \N__9872\
        );

    \I__1204\ : Span4Mux_s3_h
    port map (
            O => \N__9880\,
            I => \N__9872\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__9877\,
            I => \ufifo.fifo.rdaddrZ0Z_6\
        );

    \I__1202\ : Odrv4
    port map (
            O => \N__9872\,
            I => \ufifo.fifo.rdaddrZ0Z_6\
        );

    \I__1201\ : InMux
    port map (
            O => \N__9867\,
            I => \N__9864\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__9864\,
            I => \N__9861\
        );

    \I__1199\ : IoSpan4Mux
    port map (
            O => \N__9861\,
            I => \N__9858\
        );

    \I__1198\ : Odrv4
    port map (
            O => \N__9858\,
            I => \uart_RXD\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__9855\,
            I => \N__9849\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9854\,
            I => \N__9840\
        );

    \I__1195\ : InMux
    port map (
            O => \N__9853\,
            I => \N__9840\
        );

    \I__1194\ : InMux
    port map (
            O => \N__9852\,
            I => \N__9840\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9849\,
            I => \N__9840\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__9840\,
            I => \N__9837\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__9837\,
            I => \Lab_UT.scdp.prng_lfsr_23\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__9834\,
            I => \resetGen.N_421_cascade_\
        );

    \I__1189\ : InMux
    port map (
            O => \N__9831\,
            I => \N__9819\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9819\
        );

    \I__1187\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9819\
        );

    \I__1186\ : InMux
    port map (
            O => \N__9828\,
            I => \N__9819\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__9819\,
            I => \N__9816\
        );

    \I__1184\ : Odrv4
    port map (
            O => \N__9816\,
            I => \buart.Z_tx.N_554\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__9813\,
            I => \resetGen.N_267_cascade_\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__9810\,
            I => \N__9807\
        );

    \I__1181\ : InMux
    port map (
            O => \N__9807\,
            I => \N__9804\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__9804\,
            I => \Lab_UT.scdp.byteToEncrypt_7\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__9801\,
            I => \N__9796\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__9800\,
            I => \N__9793\
        );

    \I__1177\ : InMux
    port map (
            O => \N__9799\,
            I => \N__9783\
        );

    \I__1176\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9783\
        );

    \I__1175\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9783\
        );

    \I__1174\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9783\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__9783\,
            I => \Lab_UT.scdp.prng_lfsr_7\
        );

    \I__1172\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9768\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9768\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9778\,
            I => \N__9768\
        );

    \I__1169\ : InMux
    port map (
            O => \N__9777\,
            I => \N__9768\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__9768\,
            I => \Lab_UT.scdp.prng_lfsr_15\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__9765\,
            I => \Lab_UT.scdp.lfsrInst.N_234_i_1_cascade_\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9762\,
            I => \N__9759\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__9759\,
            I => \N__9756\
        );

    \I__1164\ : Odrv4
    port map (
            O => \N__9756\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9753\,
            I => \N__9748\
        );

    \I__1162\ : InMux
    port map (
            O => \N__9752\,
            I => \N__9745\
        );

    \I__1161\ : InMux
    port map (
            O => \N__9751\,
            I => \N__9742\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__9748\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__9745\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__9742\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9732\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__9732\,
            I => \N__9729\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__9729\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__1154\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9721\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9718\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9715\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__9721\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9718\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__9715\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9708\,
            I => \N__9702\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9699\
        );

    \I__1146\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9694\
        );

    \I__1145\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9694\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__9702\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__9699\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9694\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__9687\,
            I => \N__9684\
        );

    \I__1140\ : InMux
    port map (
            O => \N__9684\,
            I => \N__9681\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__9681\,
            I => \N__9674\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9665\
        );

    \I__1137\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9665\
        );

    \I__1136\ : InMux
    port map (
            O => \N__9678\,
            I => \N__9665\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9665\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__9674\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9665\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1132\ : IoInMux
    port map (
            O => \N__9660\,
            I => \N__9657\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__9657\,
            I => \N__9654\
        );

    \I__1130\ : Span4Mux_s1_h
    port map (
            O => \N__9654\,
            I => \N__9651\
        );

    \I__1129\ : Odrv4
    port map (
            O => \N__9651\,
            I => \buart.Z_rx.N_76_i\
        );

    \I__1128\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9645\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__9645\,
            I => \N__9642\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__9642\,
            I => \ufifo.fifo.fifo_txdata_2\
        );

    \I__1125\ : InMux
    port map (
            O => \N__9639\,
            I => \N__9636\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__9636\,
            I => \N__9633\
        );

    \I__1123\ : Odrv12
    port map (
            O => \N__9633\,
            I => \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__9630\,
            I => \ufifo.sb_ram512x8_inst_RNILSN11_cascade_\
        );

    \I__1121\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9624\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__1119\ : Odrv12
    port map (
            O => \N__9621\,
            I => utb_txdata_2
        );

    \I__1118\ : InMux
    port map (
            O => \N__9618\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__1117\ : InMux
    port map (
            O => \N__9615\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__1116\ : InMux
    port map (
            O => \N__9612\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9609\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__9606\,
            I => \N__9603\
        );

    \I__1113\ : InMux
    port map (
            O => \N__9603\,
            I => \N__9597\
        );

    \I__1112\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9597\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__9597\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__9594\,
            I => \N__9590\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9585\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9585\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__9585\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__9582\,
            I => \N__9578\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9574\
        );

    \I__1104\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9569\
        );

    \I__1103\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9569\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__9574\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__9569\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1100\ : InMux
    port map (
            O => \N__9564\,
            I => \N__9561\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__9561\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3\
        );

    \I__1098\ : InMux
    port map (
            O => \N__9558\,
            I => \N__9544\
        );

    \I__1097\ : InMux
    port map (
            O => \N__9557\,
            I => \N__9544\
        );

    \I__1096\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9544\
        );

    \I__1095\ : InMux
    port map (
            O => \N__9555\,
            I => \N__9532\
        );

    \I__1094\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9532\
        );

    \I__1093\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9532\
        );

    \I__1092\ : InMux
    port map (
            O => \N__9552\,
            I => \N__9532\
        );

    \I__1091\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9532\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__9544\,
            I => \N__9524\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9521\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__9532\,
            I => \N__9518\
        );

    \I__1087\ : InMux
    port map (
            O => \N__9531\,
            I => \N__9515\
        );

    \I__1086\ : InMux
    port map (
            O => \N__9530\,
            I => \N__9506\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9506\
        );

    \I__1084\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9506\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9506\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__9524\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__9521\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__9518\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__9515\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__9506\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__9495\,
            I => \N__9492\
        );

    \I__1076\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9479\
        );

    \I__1075\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9479\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9479\
        );

    \I__1073\ : InMux
    port map (
            O => \N__9489\,
            I => \N__9479\
        );

    \I__1072\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9474\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__9479\,
            I => \N__9471\
        );

    \I__1070\ : InMux
    port map (
            O => \N__9478\,
            I => \N__9466\
        );

    \I__1069\ : InMux
    port map (
            O => \N__9477\,
            I => \N__9466\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__9474\,
            I => \ufifo.cstate_4\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__9471\,
            I => \ufifo.cstate_4\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__9466\,
            I => \ufifo.cstate_4\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__9459\,
            I => \ufifo.tx_fsm.N_394_cascade_\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__9456\,
            I => \N__9453\
        );

    \I__1063\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9450\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__9450\,
            I => \N__9447\
        );

    \I__1061\ : Span4Mux_h
    port map (
            O => \N__9447\,
            I => \N__9442\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9446\,
            I => \N__9439\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9445\,
            I => \N__9436\
        );

    \I__1058\ : Odrv4
    port map (
            O => \N__9442\,
            I => \ufifo.fifo.wraddrZ0Z_4\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__9439\,
            I => \ufifo.fifo.wraddrZ0Z_4\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__9436\,
            I => \ufifo.fifo.wraddrZ0Z_4\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__9429\,
            I => \N__9426\
        );

    \I__1054\ : InMux
    port map (
            O => \N__9426\,
            I => \N__9423\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__9423\,
            I => \N__9419\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__9422\,
            I => \N__9415\
        );

    \I__1051\ : Span4Mux_h
    port map (
            O => \N__9419\,
            I => \N__9412\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9409\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9406\
        );

    \I__1048\ : Odrv4
    port map (
            O => \N__9412\,
            I => \ufifo.fifo.wraddrZ0Z_5\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__9409\,
            I => \ufifo.fifo.wraddrZ0Z_5\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__9406\,
            I => \ufifo.fifo.wraddrZ0Z_5\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__9399\,
            I => \N__9396\
        );

    \I__1044\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9393\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9393\,
            I => \N__9390\
        );

    \I__1042\ : Span4Mux_h
    port map (
            O => \N__9390\,
            I => \N__9385\
        );

    \I__1041\ : InMux
    port map (
            O => \N__9389\,
            I => \N__9382\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9379\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__9385\,
            I => \ufifo.fifo.wraddrZ0Z_6\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9382\,
            I => \ufifo.fifo.wraddrZ0Z_6\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__9379\,
            I => \ufifo.fifo.wraddrZ0Z_6\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__9372\,
            I => \ufifo.fifo.un1_emptyB_NE_0_cascade_\
        );

    \I__1035\ : InMux
    port map (
            O => \N__9369\,
            I => \N__9366\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__9366\,
            I => \ufifo.fifo.un1_emptyB_NE_3\
        );

    \I__1033\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9360\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__9360\,
            I => \ufifo.fifo.un1_emptyB_NE_2\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__9357\,
            I => \ufifo.fifo.un1_emptyB_NE_4_cascade_\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9354\,
            I => \N__9351\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__9351\,
            I => \ufifo.fifo.un1_emptyB_NE_1\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__9348\,
            I => \ufifo.emptyB_0_cascade_\
        );

    \I__1027\ : InMux
    port map (
            O => \N__9345\,
            I => \N__9341\
        );

    \I__1026\ : InMux
    port map (
            O => \N__9344\,
            I => \N__9338\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__9341\,
            I => \ufifo.tx_fsm.cstateZ0Z_5\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__9338\,
            I => \ufifo.tx_fsm.cstateZ0Z_5\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__9333\,
            I => \ufifo.tx_fsm.N_396_cascade_\
        );

    \I__1022\ : InMux
    port map (
            O => \N__9330\,
            I => \N__9322\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9322\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9317\
        );

    \I__1019\ : InMux
    port map (
            O => \N__9327\,
            I => \N__9317\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__9322\,
            I => \ufifo.tx_fsm.N_279\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__9317\,
            I => \ufifo.tx_fsm.N_279\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__9312\,
            I => \N__9308\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9303\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9298\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9307\,
            I => \N__9298\
        );

    \I__1012\ : InMux
    port map (
            O => \N__9306\,
            I => \N__9295\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__9303\,
            I => \ufifo.emptyB_0\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__9298\,
            I => \ufifo.emptyB_0\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__9295\,
            I => \ufifo.emptyB_0\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__9288\,
            I => \ufifo.tx_fsm.cstate_srsts_i_0_1_1_cascade_\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__9285\,
            I => \N__9280\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__9284\,
            I => \N__9277\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9274\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9271\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9268\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__9274\,
            I => \ufifo.tx_fsm.cstateZ0Z_1\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__9271\,
            I => \ufifo.tx_fsm.cstateZ0Z_1\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__9268\,
            I => \ufifo.tx_fsm.cstateZ0Z_1\
        );

    \I__999\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9258\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__9258\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__9255\,
            I => \utb_txdata_1_cascade_\
        );

    \I__996\ : InMux
    port map (
            O => \N__9252\,
            I => \N__9238\
        );

    \I__995\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9231\
        );

    \I__994\ : InMux
    port map (
            O => \N__9250\,
            I => \N__9231\
        );

    \I__993\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9231\
        );

    \I__992\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9222\
        );

    \I__991\ : InMux
    port map (
            O => \N__9247\,
            I => \N__9222\
        );

    \I__990\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9222\
        );

    \I__989\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9222\
        );

    \I__988\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9213\
        );

    \I__987\ : InMux
    port map (
            O => \N__9243\,
            I => \N__9213\
        );

    \I__986\ : InMux
    port map (
            O => \N__9242\,
            I => \N__9213\
        );

    \I__985\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9213\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__9238\,
            I => \N_257\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__9231\,
            I => \N_257\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__9222\,
            I => \N_257\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__9213\,
            I => \N_257\
        );

    \I__980\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9201\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__9201\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__978\ : CEMux
    port map (
            O => \N__9198\,
            I => \N__9193\
        );

    \I__977\ : CEMux
    port map (
            O => \N__9197\,
            I => \N__9190\
        );

    \I__976\ : CEMux
    port map (
            O => \N__9196\,
            I => \N__9187\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__9193\,
            I => \N__9184\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9190\,
            I => \N__9181\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__9187\,
            I => \N__9178\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__9184\,
            I => \buart.Z_tx.N_58\
        );

    \I__971\ : Odrv4
    port map (
            O => \N__9181\,
            I => \buart.Z_tx.N_58\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__9178\,
            I => \buart.Z_tx.N_58\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__9171\,
            I => \N__9161\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__9170\,
            I => \N__9158\
        );

    \I__967\ : InMux
    port map (
            O => \N__9169\,
            I => \N__9153\
        );

    \I__966\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9150\
        );

    \I__965\ : InMux
    port map (
            O => \N__9167\,
            I => \N__9143\
        );

    \I__964\ : InMux
    port map (
            O => \N__9166\,
            I => \N__9143\
        );

    \I__963\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9143\
        );

    \I__962\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9140\
        );

    \I__961\ : InMux
    port map (
            O => \N__9161\,
            I => \N__9131\
        );

    \I__960\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9131\
        );

    \I__959\ : InMux
    port map (
            O => \N__9157\,
            I => \N__9131\
        );

    \I__958\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9131\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__9153\,
            I => ufifo_emitcrlf_fsm_cstate_0
        );

    \I__956\ : LocalMux
    port map (
            O => \N__9150\,
            I => ufifo_emitcrlf_fsm_cstate_0
        );

    \I__955\ : LocalMux
    port map (
            O => \N__9143\,
            I => ufifo_emitcrlf_fsm_cstate_0
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9140\,
            I => ufifo_emitcrlf_fsm_cstate_0
        );

    \I__953\ : LocalMux
    port map (
            O => \N__9131\,
            I => ufifo_emitcrlf_fsm_cstate_0
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__9120\,
            I => \N__9113\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__9119\,
            I => \N__9107\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__9118\,
            I => \N__9101\
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__9117\,
            I => \N__9098\
        );

    \I__948\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9095\
        );

    \I__947\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9082\
        );

    \I__946\ : InMux
    port map (
            O => \N__9112\,
            I => \N__9082\
        );

    \I__945\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9082\
        );

    \I__944\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9082\
        );

    \I__943\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9082\
        );

    \I__942\ : InMux
    port map (
            O => \N__9106\,
            I => \N__9082\
        );

    \I__941\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9073\
        );

    \I__940\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9073\
        );

    \I__939\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9073\
        );

    \I__938\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9073\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__9095\,
            I => ufifo_emitcrlf_fsm_cstate_1
        );

    \I__936\ : LocalMux
    port map (
            O => \N__9082\,
            I => ufifo_emitcrlf_fsm_cstate_1
        );

    \I__935\ : LocalMux
    port map (
            O => \N__9073\,
            I => ufifo_emitcrlf_fsm_cstate_1
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__9066\,
            I => \N__9063\
        );

    \I__933\ : InMux
    port map (
            O => \N__9063\,
            I => \N__9060\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__9060\,
            I => \N__9057\
        );

    \I__931\ : Span4Mux_h
    port map (
            O => \N__9057\,
            I => \N__9052\
        );

    \I__930\ : InMux
    port map (
            O => \N__9056\,
            I => \N__9049\
        );

    \I__929\ : InMux
    port map (
            O => \N__9055\,
            I => \N__9046\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__9052\,
            I => \ufifo.fifo.wraddrZ0Z_2\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__9049\,
            I => \ufifo.fifo.wraddrZ0Z_2\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__9046\,
            I => \ufifo.fifo.wraddrZ0Z_2\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__9039\,
            I => \N__9036\
        );

    \I__924\ : InMux
    port map (
            O => \N__9036\,
            I => \N__9033\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__9033\,
            I => \N__9029\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__9032\,
            I => \N__9025\
        );

    \I__921\ : Span4Mux_h
    port map (
            O => \N__9029\,
            I => \N__9022\
        );

    \I__920\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9019\
        );

    \I__919\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9016\
        );

    \I__918\ : Odrv4
    port map (
            O => \N__9022\,
            I => \ufifo.fifo.wraddrZ0Z_3\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__9019\,
            I => \ufifo.fifo.wraddrZ0Z_3\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__9016\,
            I => \ufifo.fifo.wraddrZ0Z_3\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__9009\,
            I => \N__9006\
        );

    \I__914\ : InMux
    port map (
            O => \N__9006\,
            I => \N__9003\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__9003\,
            I => \N__8999\
        );

    \I__912\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8995\
        );

    \I__911\ : Span4Mux_h
    port map (
            O => \N__8999\,
            I => \N__8992\
        );

    \I__910\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8989\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__8995\,
            I => \N__8986\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__8992\,
            I => \ufifo.fifo.wraddrZ0Z_7\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__8989\,
            I => \ufifo.fifo.wraddrZ0Z_7\
        );

    \I__906\ : Odrv4
    port map (
            O => \N__8986\,
            I => \ufifo.fifo.wraddrZ0Z_7\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__8979\,
            I => \N__8975\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__8978\,
            I => \N__8972\
        );

    \I__903\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8969\
        );

    \I__902\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8966\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__8969\,
            I => \N__8960\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8960\
        );

    \I__899\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8957\
        );

    \I__898\ : Span4Mux_h
    port map (
            O => \N__8960\,
            I => \N__8954\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__8957\,
            I => \ufifo.fifo.wraddrZ0Z_8\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__8954\,
            I => \ufifo.fifo.wraddrZ0Z_8\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__8949\,
            I => \N__8946\
        );

    \I__894\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8943\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__8943\,
            I => \N__8940\
        );

    \I__892\ : Span4Mux_v
    port map (
            O => \N__8940\,
            I => \N__8935\
        );

    \I__891\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8932\
        );

    \I__890\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8929\
        );

    \I__889\ : Odrv4
    port map (
            O => \N__8935\,
            I => \ufifo.fifo.wraddrZ0Z_0\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__8932\,
            I => \ufifo.fifo.wraddrZ0Z_0\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__8929\,
            I => \ufifo.fifo.wraddrZ0Z_0\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__8922\,
            I => \N__8919\
        );

    \I__885\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8916\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__8916\,
            I => \N__8912\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__8915\,
            I => \N__8908\
        );

    \I__882\ : Span4Mux_v
    port map (
            O => \N__8912\,
            I => \N__8905\
        );

    \I__881\ : InMux
    port map (
            O => \N__8911\,
            I => \N__8902\
        );

    \I__880\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8899\
        );

    \I__879\ : Odrv4
    port map (
            O => \N__8905\,
            I => \ufifo.fifo.wraddrZ0Z_1\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__8902\,
            I => \ufifo.fifo.wraddrZ0Z_1\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__8899\,
            I => \ufifo.fifo.wraddrZ0Z_1\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__8892\,
            I => \ufifo.tx_fsm.N_358_cascade_\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__8889\,
            I => \buart.Z_tx.N_373_cascade_\
        );

    \I__874\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8883\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__8883\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__8880\,
            I => \N__8877\
        );

    \I__871\ : InMux
    port map (
            O => \N__8877\,
            I => \N__8874\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__8874\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__8871\,
            I => \N__8868\
        );

    \I__868\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8865\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__8865\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__866\ : InMux
    port map (
            O => \N__8862\,
            I => \N__8859\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__8859\,
            I => \buart.Z_tx.N_375\
        );

    \I__864\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8853\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__8853\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__8850\,
            I => \buart.Z_tx.N_215_cascade_\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__8847\,
            I => \N_257_cascade_\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__8844\,
            I => \N__8841\
        );

    \I__859\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8838\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__8838\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__8835\,
            I => \ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0_cascade_\
        );

    \I__856\ : InMux
    port map (
            O => \N__8832\,
            I => \ufifo.fifo.un1_wraddr_cry_6\
        );

    \I__855\ : InMux
    port map (
            O => \N__8829\,
            I => \bfn_1_7_0_\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__8826\,
            I => \N__8823\
        );

    \I__853\ : InMux
    port map (
            O => \N__8823\,
            I => \N__8820\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8820\,
            I => \N__8817\
        );

    \I__851\ : Span4Mux_s2_h
    port map (
            O => \N__8817\,
            I => \N__8814\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__8814\,
            I => ufifo_fifo_txdata_3
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__8811\,
            I => \buart.Z_tx.N_369_cascade_\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__8808\,
            I => \N__8805\
        );

    \I__847\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8802\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__8802\,
            I => \N__8799\
        );

    \I__845\ : Span4Mux_s2_h
    port map (
            O => \N__8799\,
            I => \N__8796\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__8796\,
            I => ufifo_fifo_txdata_4
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__8793\,
            I => \buart.Z_tx.N_371_cascade_\
        );

    \I__842\ : InMux
    port map (
            O => \N__8790\,
            I => \N__8787\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__8787\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__840\ : InMux
    port map (
            O => \N__8784\,
            I => \N__8774\
        );

    \I__839\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8774\
        );

    \I__838\ : InMux
    port map (
            O => \N__8782\,
            I => \N__8774\
        );

    \I__837\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8771\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8774\,
            I => \N_366\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__8771\,
            I => \N_366\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__8766\,
            I => \N__8763\
        );

    \I__833\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8760\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__8760\,
            I => \N__8757\
        );

    \I__831\ : Span4Mux_s2_v
    port map (
            O => \N__8757\,
            I => \N__8754\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__8754\,
            I => ufifo_fifo_txdata_5
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__8751\,
            I => \ufifo.emitcrlf_fsm.N_501_cascade_\
        );

    \I__828\ : InMux
    port map (
            O => \N__8748\,
            I => \N__8745\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__8745\,
            I => \ufifo.emitcrlf_fsm.cstate_ns_i_0_0_1\
        );

    \I__826\ : InMux
    port map (
            O => \N__8742\,
            I => \ufifo.fifo.un1_wraddr_cry_0\
        );

    \I__825\ : InMux
    port map (
            O => \N__8739\,
            I => \ufifo.fifo.un1_wraddr_cry_1\
        );

    \I__824\ : InMux
    port map (
            O => \N__8736\,
            I => \ufifo.fifo.un1_wraddr_cry_2\
        );

    \I__823\ : InMux
    port map (
            O => \N__8733\,
            I => \ufifo.fifo.un1_wraddr_cry_3\
        );

    \I__822\ : InMux
    port map (
            O => \N__8730\,
            I => \ufifo.fifo.un1_wraddr_cry_4\
        );

    \I__821\ : InMux
    port map (
            O => \N__8727\,
            I => \ufifo.fifo.un1_wraddr_cry_5\
        );

    \I__820\ : InMux
    port map (
            O => \N__8724\,
            I => \N__8721\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__8721\,
            I => \N__8718\
        );

    \I__818\ : Span4Mux_s2_h
    port map (
            O => \N__8718\,
            I => \N__8715\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__8715\,
            I => \ufifo.fifo.fifo_txdata_7\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__8712\,
            I => \N_366_cascade_\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__8709\,
            I => \ufifo_utb_txdata_m0_7_cascade_\
        );

    \I__814\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8703\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__8703\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__8700\,
            I => \ufifo.emitcrlf_fsm.cstate_ns_i_0_2_1_cascade_\
        );

    \I__811\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8694\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__8694\,
            I => \ufifo.N_323\
        );

    \I__809\ : CascadeMux
    port map (
            O => \N__8691\,
            I => \buart.Z_tx.un1_bitcount_c3_cascade_\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__8688\,
            I => \N__8684\
        );

    \I__807\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8679\
        );

    \I__806\ : InMux
    port map (
            O => \N__8684\,
            I => \N__8679\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__8679\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__8676\,
            I => \ufifo_utb_txdata_rdy_0_i_1_cascade_\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__8673\,
            I => \N__8668\
        );

    \I__802\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8664\
        );

    \I__801\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8657\
        );

    \I__800\ : InMux
    port map (
            O => \N__8668\,
            I => \N__8657\
        );

    \I__799\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8657\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__8664\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8657\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__796\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8645\
        );

    \I__795\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8636\
        );

    \I__794\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8636\
        );

    \I__793\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8636\
        );

    \I__792\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8636\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__8645\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__8636\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__789\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8628\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__8628\,
            I => \buart.Z_tx.un1_bitcount_c2\
        );

    \I__787\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8619\
        );

    \I__786\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8619\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__8619\,
            I => ufifo_utb_txdata_rdy_0_i_1
        );

    \I__784\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8607\
        );

    \I__783\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8607\
        );

    \I__782\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8607\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__8607\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__8604\,
            I => \N__8599\
        );

    \I__779\ : InMux
    port map (
            O => \N__8603\,
            I => \N__8591\
        );

    \I__778\ : InMux
    port map (
            O => \N__8602\,
            I => \N__8591\
        );

    \I__777\ : InMux
    port map (
            O => \N__8599\,
            I => \N__8582\
        );

    \I__776\ : InMux
    port map (
            O => \N__8598\,
            I => \N__8582\
        );

    \I__775\ : InMux
    port map (
            O => \N__8597\,
            I => \N__8582\
        );

    \I__774\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8582\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__8591\,
            I => \buart.Z_tx.counter_RNIVE1P1_0\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8582\,
            I => \buart.Z_tx.counter_RNIVE1P1_0\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__8577\,
            I => \N__8574\
        );

    \I__770\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8571\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__8571\,
            I => \N__8568\
        );

    \I__768\ : Span4Mux_s2_h
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__767\ : Odrv4
    port map (
            O => \N__8565\,
            I => ufifo_fifo_txdata_6
        );

    \I__766\ : IoInMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__8559\,
            I => \N__8556\
        );

    \I__764\ : IoSpan4Mux
    port map (
            O => \N__8556\,
            I => \N__8553\
        );

    \I__763\ : IoSpan4Mux
    port map (
            O => \N__8553\,
            I => \N__8550\
        );

    \I__762\ : Odrv4
    port map (
            O => \N__8550\,
            I => o_serial_data_c
        );

    \I__761\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8544\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__8544\,
            I => \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_6\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__8541\,
            I => \N__8537\
        );

    \I__758\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8532\
        );

    \I__757\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8532\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__8532\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__8529\,
            I => \N__8526\
        );

    \I__754\ : InMux
    port map (
            O => \N__8526\,
            I => \N__8523\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__8523\,
            I => \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_5\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__8520\,
            I => \N__8517\
        );

    \I__751\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8511\
        );

    \I__750\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8511\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__8511\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__748\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8504\
        );

    \I__747\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8501\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__8504\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8501\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__744\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8491\
        );

    \I__743\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8486\
        );

    \I__742\ : InMux
    port map (
            O => \N__8494\,
            I => \N__8486\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__8491\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__8486\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__8481\,
            I => \N__8477\
        );

    \I__738\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8473\
        );

    \I__737\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8468\
        );

    \I__736\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8468\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__8473\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_0\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__8468\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_0\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__8463\,
            I => \N__8459\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__8462\,
            I => \N__8451\
        );

    \I__731\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8440\
        );

    \I__730\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8440\
        );

    \I__729\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8440\
        );

    \I__728\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8440\
        );

    \I__727\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8440\
        );

    \I__726\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8435\
        );

    \I__725\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8435\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__8440\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__8435\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__722\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8421\
        );

    \I__721\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8421\
        );

    \I__720\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8421\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__8421\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__8418\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_0_cascade_\
        );

    \I__717\ : CascadeMux
    port map (
            O => \N__8415\,
            I => \buart.Z_tx.counter_RNIVE1P1_0_cascade_\
        );

    \I__716\ : InMux
    port map (
            O => \N__8412\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__715\ : InMux
    port map (
            O => \N__8409\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__714\ : InMux
    port map (
            O => \N__8406\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__713\ : InMux
    port map (
            O => \N__8403\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__712\ : InMux
    port map (
            O => \N__8400\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__8397\,
            I => \N__8394\
        );

    \I__710\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8388\
        );

    \I__709\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8388\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__8388\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__707\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8382\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__8382\,
            I => \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_3\
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__8379\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_\
        );

    \I__704\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8370\
        );

    \I__703\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8370\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__8370\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__701\ : IoInMux
    port map (
            O => \N__8367\,
            I => \N__8364\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__8364\,
            I => \N__8361\
        );

    \I__699\ : Span12Mux_s9_v
    port map (
            O => \N__8361\,
            I => \N__8358\
        );

    \I__698\ : Odrv12
    port map (
            O => \N__8358\,
            I => \latticehx1k_pll_inst.clk\
        );

    \I__697\ : IoInMux
    port map (
            O => \N__8355\,
            I => \N__8352\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__8352\,
            I => \N__8349\
        );

    \I__695\ : IoSpan4Mux
    port map (
            O => \N__8349\,
            I => \N__8346\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__8346\,
            I => clk_in_c
        );

    \IN_MUX_bfv_1_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_1_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ufifo.fifo.un1_wraddr_cry_7\,
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_4_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_4_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ufifo.fifo.un1_rdaddr_cry_7\,
            carryinitout => \bfn_4_5_0_\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8367\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \resetGen.rst_1_iso_RNIU3O8\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__16451\,
            GLOBALBUFFEROUTPUT => \resetGen_rst_1_iso_g\
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9660\,
            GLOBALBUFFEROUTPUT => \N_76_i_g\
        );

    \Lab_UT.scctrl.state_1_ret_5_RNI\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10530\,
            GLOBALBUFFEROUTPUT => \Lab_UT.sccLdLFSR_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8496\,
            in2 => \N__8462\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_1_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8397\,
            in3 => \N__8412\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__21150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNO_0_3_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8376\,
            in2 => \_gnd_net_\,
            in3 => \N__8409\,
            lcout => \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8508\,
            in2 => \_gnd_net_\,
            in3 => \N__8406\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__21150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNO_0_5_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8520\,
            in3 => \N__8403\,
            lcout => \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNO_0_6_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8540\,
            in2 => \_gnd_net_\,
            in3 => \N__8400\,
            lcout => \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIGU38_6_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8516\,
            in1 => \N__8375\,
            in2 => \N__8541\,
            in3 => \N__8393\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__8480\,
            in1 => \N__8385\,
            in2 => \N__8379\,
            in3 => \N__8454\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__8458\,
            in1 => \N__8547\,
            in2 => \N__8481\,
            in3 => \N__8430\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__8429\,
            in1 => \N__8476\,
            in2 => \N__8529\,
            in3 => \N__8457\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8456\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__8495\,
            in1 => \_gnd_net_\,
            in2 => \N__8463\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21149\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5S14_1_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8507\,
            in2 => \_gnd_net_\,
            in3 => \N__8494\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_0\,
            ltout => \buart.Z_tx.Z_baudgen.ser_clk_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_0_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8455\,
            in1 => \N__8428\,
            in2 => \N__8418\,
            in3 => \N__9543\,
            lcout => \buart.Z_tx.counter_RNIVE1P1_0\,
            ltout => \buart.Z_tx.counter_RNIVE1P1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8672\,
            in2 => \N__8415\,
            in3 => \N__8652\,
            lcout => \buart.Z_tx.un1_bitcount_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIQOQA1_3_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8614\,
            in1 => \N__8667\,
            in2 => \N__8688\,
            in3 => \N__8648\,
            lcout => \buart__tx_uart_busy_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__8649\,
            in1 => \N__8596\,
            in2 => \N__8673\,
            in3 => \N__8615\,
            lcout => OPEN,
            ltout => \buart.Z_tx.un1_bitcount_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_3_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110010110"
        )
    port map (
            in0 => \N__8687\,
            in1 => \N__8603\,
            in2 => \N__8691\,
            in3 => \N__8625\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21148\,
            ce => 'H',
            sr => \N__20833\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIPKRF7_0_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12320\,
            in2 => \_gnd_net_\,
            in3 => \N__9249\,
            lcout => ufifo_utb_txdata_rdy_0_i_1,
            ltout => \ufifo_utb_txdata_rdy_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_1_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011110110"
        )
    port map (
            in0 => \N__8598\,
            in1 => \N__8671\,
            in2 => \N__8676\,
            in3 => \N__8650\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21148\,
            ce => 'H',
            sr => \N__20833\
        );

    \buart.Z_tx.bitcount_0_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8651\,
            in1 => \N__8597\,
            in2 => \_gnd_net_\,
            in3 => \N__9251\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21148\,
            ce => 'H',
            sr => \N__20833\
        );

    \buart.Z_tx.bitcount_2_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010010110"
        )
    port map (
            in0 => \N__8616\,
            in1 => \N__8631\,
            in2 => \N__8604\,
            in3 => \N__8624\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21148\,
            ce => 'H',
            sr => \N__20833\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIO3T89_0_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__8602\,
            in1 => \N__12321\,
            in2 => \_gnd_net_\,
            in3 => \N__9250\,
            lcout => \buart.Z_tx.N_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_RNO_0_7_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__8781\,
            in1 => \N__14935\,
            in2 => \N__8577\,
            in3 => \N__9241\,
            lcout => \buart.Z_tx.N_375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.uart_tx_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9244\,
            in1 => \N__8706\,
            in2 => \_gnd_net_\,
            in3 => \N__12315\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21146\,
            ce => \N__9196\,
            sr => \N__20831\
        );

    \ufifo.tx_fsm.cstate_RNI57IK1_0_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__9168\,
            in1 => \N__9116\,
            in2 => \N__10412\,
            in3 => \N__9531\,
            lcout => \N_366\,
            ltout => \N_366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNIEQME2_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8724\,
            in2 => \N__8712\,
            in3 => \N__14529\,
            lcout => OPEN,
            ltout => \ufifo_utb_txdata_m0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_8_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001010101"
        )
    port map (
            in0 => \N__12314\,
            in1 => \_gnd_net_\,
            in2 => \N__8709\,
            in3 => \N__9243\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21146\,
            ce => \N__9196\,
            sr => \N__20831\
        );

    \buart.Z_tx.shifter_0_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__9242\,
            in1 => \_gnd_net_\,
            in2 => \N__8844\,
            in3 => \N__12313\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21146\,
            ce => \N__9196\,
            sr => \N__20831\
        );

    \ufifo.emitcrlf_fsm.cstate_RNO_0_1_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100100"
        )
    port map (
            in0 => \N__9554\,
            in1 => \N__9111\,
            in2 => \N__9171\,
            in3 => \N__8748\,
            lcout => OPEN,
            ltout => \ufifo.emitcrlf_fsm.cstate_ns_i_0_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_1_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__9112\,
            in1 => \N__8697\,
            in2 => \N__8700\,
            in3 => \N__15449\,
            lcout => ufifo_emitcrlf_fsm_cstate_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21144\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNI7ELR5_4_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__9553\,
            in1 => \N__9478\,
            in2 => \_gnd_net_\,
            in3 => \N__9306\,
            lcout => \ufifo.N_323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_0_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101000000000"
        )
    port map (
            in0 => \N__9169\,
            in1 => \N__9555\,
            in2 => \N__9120\,
            in3 => \N__15448\,
            lcout => ufifo_emitcrlf_fsm_cstate_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21144\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_srsts_i_i_o2_2_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101111111"
        )
    port map (
            in0 => \N__9552\,
            in1 => \N__9110\,
            in2 => \N__9170\,
            in3 => \_gnd_net_\,
            lcout => \ufifo.tx_fsm.N_279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_0_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9551\,
            in2 => \N__9119\,
            in3 => \N__9156\,
            lcout => \N_368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNO_2_1_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__9157\,
            in1 => \N__9106\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \ufifo.emitcrlf_fsm.N_501_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNO_1_1_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__9477\,
            in1 => \N__10401\,
            in2 => \N__8751\,
            in3 => \N__23208\,
            lcout => \ufifo.emitcrlf_fsm.cstate_ns_i_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_0_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8939\,
            in2 => \N__11303\,
            in3 => \N__11301\,
            lcout => \ufifo.fifo.wraddrZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \ufifo.fifo.un1_wraddr_cry_0\,
            clk => \N__21140\,
            ce => 'H',
            sr => \N__20808\
        );

    \ufifo.fifo.wraddr_1_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8911\,
            in2 => \_gnd_net_\,
            in3 => \N__8742\,
            lcout => \ufifo.fifo.wraddrZ0Z_1\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_0\,
            carryout => \ufifo.fifo.un1_wraddr_cry_1\,
            clk => \N__21140\,
            ce => 'H',
            sr => \N__20808\
        );

    \ufifo.fifo.wraddr_2_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9056\,
            in2 => \_gnd_net_\,
            in3 => \N__8739\,
            lcout => \ufifo.fifo.wraddrZ0Z_2\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_1\,
            carryout => \ufifo.fifo.un1_wraddr_cry_2\,
            clk => \N__21140\,
            ce => 'H',
            sr => \N__20808\
        );

    \ufifo.fifo.wraddr_3_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9028\,
            in2 => \_gnd_net_\,
            in3 => \N__8736\,
            lcout => \ufifo.fifo.wraddrZ0Z_3\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_2\,
            carryout => \ufifo.fifo.un1_wraddr_cry_3\,
            clk => \N__21140\,
            ce => 'H',
            sr => \N__20808\
        );

    \ufifo.fifo.wraddr_4_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9446\,
            in2 => \_gnd_net_\,
            in3 => \N__8733\,
            lcout => \ufifo.fifo.wraddrZ0Z_4\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_3\,
            carryout => \ufifo.fifo.un1_wraddr_cry_4\,
            clk => \N__21140\,
            ce => 'H',
            sr => \N__20808\
        );

    \ufifo.fifo.wraddr_5_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9418\,
            in2 => \_gnd_net_\,
            in3 => \N__8730\,
            lcout => \ufifo.fifo.wraddrZ0Z_5\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_4\,
            carryout => \ufifo.fifo.un1_wraddr_cry_5\,
            clk => \N__21140\,
            ce => 'H',
            sr => \N__20808\
        );

    \ufifo.fifo.wraddr_6_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9389\,
            in2 => \_gnd_net_\,
            in3 => \N__8727\,
            lcout => \ufifo.fifo.wraddrZ0Z_6\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_5\,
            carryout => \ufifo.fifo.un1_wraddr_cry_6\,
            clk => \N__21140\,
            ce => 'H',
            sr => \N__20808\
        );

    \ufifo.fifo.wraddr_7_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8998\,
            in2 => \_gnd_net_\,
            in3 => \N__8832\,
            lcout => \ufifo.fifo.wraddrZ0Z_7\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_6\,
            carryout => \ufifo.fifo.un1_wraddr_cry_7\,
            clk => \N__21140\,
            ce => 'H',
            sr => \N__20808\
        );

    \ufifo.fifo.wraddr_8_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8965\,
            in2 => \_gnd_net_\,
            in3 => \N__8829\,
            lcout => \ufifo.fifo.wraddrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21132\,
            ce => 'H',
            sr => \N__20807\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__9705\,
            in1 => \N__9724\,
            in2 => \_gnd_net_\,
            in3 => \N__9564\,
            lcout => \buart.Z_rx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__9581\,
            in1 => \N__17703\,
            in2 => \_gnd_net_\,
            in3 => \N__9706\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.EmsBitsSl_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10827\,
            lcout => \Lab_UT.sccEmsBitsSl\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21108\,
            ce => 'H',
            sr => \N__20810\
        );

    \buart.Z_tx.shifter_RNO_0_4_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__8782\,
            in1 => \N__13551\,
            in2 => \N__8826\,
            in3 => \N__9245\,
            lcout => OPEN,
            ltout => \buart.Z_tx.N_369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_4_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__12322\,
            in1 => \N__8790\,
            in2 => \N__8811\,
            in3 => \N__9828\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__9197\,
            sr => \N__20838\
        );

    \buart.Z_tx.shifter_RNO_0_5_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001001100"
        )
    port map (
            in0 => \N__8783\,
            in1 => \N__9246\,
            in2 => \N__8808\,
            in3 => \N__15127\,
            lcout => OPEN,
            ltout => \buart.Z_tx.N_371_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_5_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__12323\,
            in1 => \N__8886\,
            in2 => \N__8793\,
            in3 => \N__9829\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__9197\,
            sr => \N__20838\
        );

    \buart.Z_tx.shifter_RNO_0_6_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001001100"
        )
    port map (
            in0 => \N__8784\,
            in1 => \N__9247\,
            in2 => \N__8766\,
            in3 => \N__18808\,
            lcout => OPEN,
            ltout => \buart.Z_tx.N_373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_6_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__12324\,
            in1 => \N__8856\,
            in2 => \N__8889\,
            in3 => \N__9830\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__9197\,
            sr => \N__20838\
        );

    \buart.Z_tx.shifter_3_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__9627\,
            in1 => \N__12326\,
            in2 => \N__8880\,
            in3 => \N__9248\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__9197\,
            sr => \N__20838\
        );

    \buart.Z_tx.shifter_7_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__12325\,
            in1 => \N__9831\,
            in2 => \N__8871\,
            in3 => \N__8862\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21147\,
            ce => \N__9197\,
            sr => \N__20838\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2_0_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9529\,
            in1 => \N__9104\,
            in2 => \_gnd_net_\,
            in3 => \N__9165\,
            lcout => \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIF2CB3_3_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100011111111"
        )
    port map (
            in0 => \N__9166\,
            in1 => \N__9527\,
            in2 => \N__9117\,
            in3 => \N__14383\,
            lcout => OPEN,
            ltout => \buart.Z_tx.N_215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNI6VV36_3_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110110011"
        )
    port map (
            in0 => \N__11121\,
            in1 => \N__10205\,
            in2 => \N__8850\,
            in3 => \N__10269\,
            lcout => \N_257\,
            ltout => \N_257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__9204\,
            in1 => \N__12255\,
            in2 => \N__8847\,
            in3 => \N__12311\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21145\,
            ce => \N__9198\,
            sr => \N__20835\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__9530\,
            in1 => \N__9105\,
            in2 => \_gnd_net_\,
            in3 => \N__9167\,
            lcout => OPEN,
            ltout => \ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIQ6FP3_0_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10239\,
            in2 => \N__8835\,
            in3 => \N__12310\,
            lcout => OPEN,
            ltout => \utb_txdata_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_2_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__12312\,
            in1 => \N__9261\,
            in2 => \N__9255\,
            in3 => \N__9252\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21145\,
            ce => \N__9198\,
            sr => \N__20835\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1_0_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9164\,
            in2 => \N__9118\,
            in3 => \N__9528\,
            lcout => \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_RNIOP7U_2_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__9055\,
            in1 => \N__9986\,
            in2 => \N__9032\,
            in3 => \N__10022\,
            lcout => \ufifo.fifo.un1_emptyB_NE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_RNICE8U_8_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__9002\,
            in1 => \N__10292\,
            in2 => \N__8978\,
            in3 => \N__10322\,
            lcout => \ufifo.fifo.un1_emptyB_NE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_RNIGH7U_0_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__8938\,
            in1 => \N__10049\,
            in2 => \N__8915\,
            in3 => \N__10085\,
            lcout => \ufifo.fifo.un1_emptyB_NE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNO_0_2_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__9490\,
            in1 => \N__9307\,
            in2 => \N__9284\,
            in3 => \N__9556\,
            lcout => OPEN,
            ltout => \ufifo.tx_fsm.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_2_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__20176\,
            in1 => \N__9491\,
            in2 => \N__8892\,
            in3 => \N__9329\,
            lcout => \ufifo.popFifo\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_4_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110010"
        )
    port map (
            in0 => \N__10227\,
            in1 => \N__20177\,
            in2 => \N__9495\,
            in3 => \N__9558\,
            lcout => \ufifo.cstate_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNO_0_5_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__9557\,
            in1 => \N__9344\,
            in2 => \N__9312\,
            in3 => \N__9489\,
            lcout => OPEN,
            ltout => \ufifo.tx_fsm.N_394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_5_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__9330\,
            in1 => \N__9488\,
            in2 => \N__9459\,
            in3 => \N__20178\,
            lcout => \ufifo.tx_fsm.cstateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_RNI028U_4_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__9445\,
            in1 => \N__9926\,
            in2 => \N__9422\,
            in3 => \N__9953\,
            lcout => OPEN,
            ltout => \ufifo.fifo.un1_emptyB_NE_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_RNI36CD1_6_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9388\,
            in2 => \N__9372\,
            in3 => \N__9893\,
            lcout => OPEN,
            ltout => \ufifo.fifo.un1_emptyB_NE_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_RNINV384_0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9369\,
            in1 => \N__9363\,
            in2 => \N__9357\,
            in3 => \N__9354\,
            lcout => \ufifo.emptyB_0\,
            ltout => \ufifo.emptyB_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNO_0_0_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10402\,
            in2 => \N__9348\,
            in3 => \N__23210\,
            lcout => OPEN,
            ltout => \ufifo.tx_fsm.N_396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstateZ0Z_0_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__20175\,
            in1 => \N__9345\,
            in2 => \N__9333\,
            in3 => \N__9328\,
            lcout => ufifo_tx_fsm_cstate_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNO_0_1_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011100"
        )
    port map (
            in0 => \N__9327\,
            in1 => \N__10403\,
            in2 => \N__9285\,
            in3 => \N__23211\,
            lcout => OPEN,
            ltout => \ufifo.tx_fsm.cstate_srsts_i_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_1_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101000000000"
        )
    port map (
            in0 => \N__9283\,
            in1 => \N__9311\,
            in2 => \N__9288\,
            in3 => \N__15459\,
            lcout => \ufifo.tx_fsm.cstateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNILSN11_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9648\,
            in1 => \N__10400\,
            in2 => \_gnd_net_\,
            in3 => \N__13032\,
            lcout => OPEN,
            ltout => \ufifo.sb_ram512x8_inst_RNILSN11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIR7FP3_0_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9639\,
            in2 => \N__9630\,
            in3 => \N__12316\,
            lcout => utb_txdata_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9707\,
            in2 => \N__9582\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9725\,
            in2 => \_gnd_net_\,
            in3 => \N__9618\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__17702\,
            in1 => \_gnd_net_\,
            in2 => \N__9606\,
            in3 => \N__9615\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__21116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9752\,
            in2 => \_gnd_net_\,
            in3 => \N__9612\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__17701\,
            in1 => \N__9593\,
            in2 => \N__9687\,
            in3 => \N__9609\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9751\,
            in1 => \N__9602\,
            in2 => \N__9594\,
            in3 => \N__9577\,
            lcout => \buart.Z_rx.Z_baudgen.ser_clk_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__9680\,
            in1 => \N__9762\,
            in2 => \N__17700\,
            in3 => \N__9753\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__9679\,
            in1 => \N__9735\,
            in2 => \N__17699\,
            in3 => \N__9726\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9708\,
            in2 => \_gnd_net_\,
            in3 => \N__17685\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIELQA6_0_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__9678\,
            in1 => \N__17793\,
            in2 => \N__17698\,
            in3 => \N__14366\,
            lcout => \buart.Z_rx.N_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__11324\,
            in1 => \N__9677\,
            in2 => \N__11340\,
            in3 => \N__13869\,
            lcout => \buart.Z_rx.N_76_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u2.q_esr_0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16580\,
            lcout => \Lab_UT.scdp.byteToEncrypt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21100\,
            ce => \N__13905\,
            sr => \N__20811\
        );

    \Lab_UT.scdp.u2.q_esr_1_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17205\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scdp.byteToEncrypt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21100\,
            ce => \N__13905\,
            sr => \N__20811\
        );

    \Lab_UT.scdp.u2.q_esr_2_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13033\,
            lcout => \Lab_UT.scdp.byteToEncrypt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21100\,
            ce => \N__13905\,
            sr => \N__20811\
        );

    \Lab_UT.scdp.u2.q_esr_3_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13548\,
            lcout => \Lab_UT.scdp.byteToEncrypt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21100\,
            ce => \N__13905\,
            sr => \N__20811\
        );

    \Lab_UT.scdp.u2.q_esr_4_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15128\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scdp.byteToEncrypt_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21100\,
            ce => \N__13905\,
            sr => \N__20811\
        );

    \Lab_UT.scdp.u2.q_esr_5_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18813\,
            lcout => \Lab_UT.scdp.byteToEncrypt_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21100\,
            ce => \N__13905\,
            sr => \N__20811\
        );

    \Lab_UT.scdp.u2.q_esr_6_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14940\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scdp.byteToEncrypt_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21100\,
            ce => \N__13905\,
            sr => \N__20811\
        );

    \Lab_UT.scdp.u2.q_esr_7_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14528\,
            lcout => \Lab_UT.scdp.byteToEncrypt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21100\,
            ce => \N__13905\,
            sr => \N__20811\
        );

    \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_3_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9799\,
            in1 => \N__9854\,
            in2 => \N__9810\,
            in3 => \N__9780\,
            lcout => \Lab_UT.scdp.b2a0.N_227_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_1_7_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16928\,
            in1 => \N__9852\,
            in2 => \N__9800\,
            in3 => \N__9778\,
            lcout => \Lab_UT.scdp.lfsrInst.N_234_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_7_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9777\,
            in1 => \N__9792\,
            in2 => \N__9855\,
            in3 => \N__16927\,
            lcout => \Lab_UT.scdp.N_234_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_7_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11436\,
            lcout => \Lab_UT.scdp.prng_lfsr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21095\,
            ce => \N__12792\,
            sr => \N__20834\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_15_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14154\,
            lcout => \Lab_UT.scdp.prng_lfsr_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21095\,
            ce => \N__12792\,
            sr => \N__20834\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_0_7_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16929\,
            in1 => \N__9853\,
            in2 => \N__9801\,
            in3 => \N__9779\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.lfsrInst.N_234_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNILRI45_7_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101111111"
        )
    port map (
            in0 => \N__11460\,
            in1 => \N__11583\,
            in2 => \N__9765\,
            in3 => \N__11553\,
            lcout => \Lab_UT.scdp.g0_0_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_0_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9867\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21090\,
            ce => 'H',
            sr => \N__20837\
        );

    \buart.Z_rx.hh_1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17762\,
            lcout => \buart__rx_hh_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21090\,
            ce => 'H',
            sr => \N__20837\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_23_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18459\,
            lcout => \Lab_UT.scdp.prng_lfsr_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21084\,
            ce => \N__12791\,
            sr => \N__20841\
        );

    \resetGen.shifter_ret_RNIC2S44_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10267\,
            in1 => \N__15125\,
            in2 => \_gnd_net_\,
            in3 => \N__14381\,
            lcout => \resetGen.N_421\,
            ltout => \resetGen.N_421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__22561\,
            in1 => \_gnd_net_\,
            in2 => \N__9834\,
            in3 => \N__10181\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_4_0_o2_2_4_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__10268\,
            in1 => \N__15126\,
            in2 => \N__10206\,
            in3 => \N__14382\,
            lcout => \buart.Z_tx.N_554\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010110100"
        )
    port map (
            in0 => \N__22562\,
            in1 => \N__10182\,
            in2 => \N__10167\,
            in3 => \N__10444\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNO_0_2_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__10180\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10163\,
            lcout => OPEN,
            ltout => \resetGen.N_267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001001"
        )
    port map (
            in0 => \N__22563\,
            in1 => \N__10152\,
            in2 => \N__9813\,
            in3 => \N__10445\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNITEEC1_2_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__10179\,
            in1 => \N__10162\,
            in2 => \_gnd_net_\,
            in3 => \N__10151\,
            lcout => \resetGen.N_274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_3_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10135\,
            in2 => \_gnd_net_\,
            in3 => \N__15458\,
            lcout => ufifo_fifo_txdata_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.rdaddr_0_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10075\,
            in2 => \N__10139\,
            in3 => \N__10134\,
            lcout => \ufifo.fifo.rdaddrZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_4_0_\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_0\,
            clk => \N__21136\,
            ce => 'H',
            sr => \N__20818\
        );

    \ufifo.fifo.rdaddr_1_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10042\,
            in2 => \_gnd_net_\,
            in3 => \N__10026\,
            lcout => \ufifo.fifo.rdaddrZ0Z_1\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_0\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_1\,
            clk => \N__21136\,
            ce => 'H',
            sr => \N__20818\
        );

    \ufifo.fifo.rdaddr_2_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10012\,
            in2 => \_gnd_net_\,
            in3 => \N__9993\,
            lcout => \ufifo.fifo.rdaddrZ0Z_2\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_1\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_2\,
            clk => \N__21136\,
            ce => 'H',
            sr => \N__20818\
        );

    \ufifo.fifo.rdaddr_3_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9979\,
            in2 => \_gnd_net_\,
            in3 => \N__9960\,
            lcout => \ufifo.fifo.rdaddrZ0Z_3\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_2\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_3\,
            clk => \N__21136\,
            ce => 'H',
            sr => \N__20818\
        );

    \ufifo.fifo.rdaddr_4_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9946\,
            in2 => \_gnd_net_\,
            in3 => \N__9930\,
            lcout => \ufifo.fifo.rdaddrZ0Z_4\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_3\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_4\,
            clk => \N__21136\,
            ce => 'H',
            sr => \N__20818\
        );

    \ufifo.fifo.rdaddr_5_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9919\,
            in2 => \_gnd_net_\,
            in3 => \N__9900\,
            lcout => \ufifo.fifo.rdaddrZ0Z_5\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_4\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_5\,
            clk => \N__21136\,
            ce => 'H',
            sr => \N__20818\
        );

    \ufifo.fifo.rdaddr_6_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9886\,
            in2 => \_gnd_net_\,
            in3 => \N__10329\,
            lcout => \ufifo.fifo.rdaddrZ0Z_6\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_5\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_6\,
            clk => \N__21136\,
            ce => 'H',
            sr => \N__20818\
        );

    \ufifo.fifo.rdaddr_7_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10321\,
            in2 => \_gnd_net_\,
            in3 => \N__10299\,
            lcout => \ufifo.fifo.rdaddrZ0Z_7\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_6\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_7\,
            clk => \N__21136\,
            ce => 'H',
            sr => \N__20818\
        );

    \ufifo.fifo.rdaddr_8_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10288\,
            in2 => \_gnd_net_\,
            in3 => \N__10296\,
            lcout => \ufifo.fifo.rdaddrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21127\,
            ce => 'H',
            sr => \N__20815\
        );

    \resetGen.shifter_ret_RNITHBO1_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__13010\,
            in1 => \N__11130\,
            in2 => \N__17190\,
            in3 => \N__17022\,
            lcout => \N_251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_esr_2_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__17023\,
            in1 => \N__17160\,
            in2 => \N__13038\,
            in3 => \N__16642\,
            lcout => \Lab_UT.scdp.u0.byteToDecrypt_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21122\,
            ce => \N__16410\,
            sr => \N__20814\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNIKRN11_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10245\,
            in1 => \N__10405\,
            in2 => \_gnd_net_\,
            in3 => \N__17159\,
            lcout => \ufifo.sb_ram512x8_inst_RNIKRN11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_4_0_o2_3_4_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__10404\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10223\,
            lcout => \buart.Z_tx.N_278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__22539\,
            in1 => \N__10464\,
            in2 => \N__10431\,
            in3 => \N__10452\,
            lcout => rst_ii,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.state_1_ret_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22541\,
            lcout => rst_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100001"
        )
    port map (
            in0 => \N__22538\,
            in1 => \N__10463\,
            in2 => \N__10430\,
            in3 => \N__10451\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNIKTQ21_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10416\,
            in1 => \N__10356\,
            in2 => \_gnd_net_\,
            in3 => \N__16562\,
            lcout => \ufifo.sb_ram512x8_inst_RNIKTQ21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_1_iso_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22540\,
            lcout => \resetGen_rst_1_iso\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_3_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17735\,
            in2 => \_gnd_net_\,
            in3 => \N__14909\,
            lcout => \N_233_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNI679E_6_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10665\,
            in1 => \N__10491\,
            in2 => \_gnd_net_\,
            in3 => \N__10836\,
            lcout => \Lab_UT.scdp.msBitsi.q_esr_RNI679EZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lsBitsi.q_esr_2_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__10539\,
            in1 => \N__10556\,
            in2 => \N__10590\,
            in3 => \N__12638\,
            lcout => \Lab_UT.scdp.lsBitsD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21110\,
            ce => \N__11217\,
            sr => \N__20809\
        );

    \Lab_UT.scdp.lsBitsi.q_esr_4_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100111111111"
        )
    port map (
            in0 => \N__12639\,
            in1 => \N__10588\,
            in2 => \N__10560\,
            in3 => \N__11693\,
            lcout => \Lab_UT.scdp.lsBitsD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21110\,
            ce => \N__11217\,
            sr => \N__20809\
        );

    \Lab_UT.scdp.b2a1.asciiHex_2_i_o2_2_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__11691\,
            in1 => \N__10343\,
            in2 => \_gnd_net_\,
            in3 => \N__12707\,
            lcout => \Lab_UT.scdp.b2a1.N_293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lsBitsi.q_esr_0_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__12708\,
            in1 => \N__10476\,
            in2 => \N__10347\,
            in3 => \N__11692\,
            lcout => \Lab_UT.scdp.lsBitsD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21110\,
            ce => \N__11217\,
            sr => \N__20809\
        );

    \Lab_UT.scdp.b2a1.lsBits_i_0_o2_6_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010101010111"
        )
    port map (
            in0 => \N__11690\,
            in1 => \N__10554\,
            in2 => \N__10589\,
            in3 => \N__12636\,
            lcout => \Lab_UT.scdp.lsBits_i_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.b2a1.asciiHex_2_i_x2_0_2_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10602\,
            in1 => \N__11847\,
            in2 => \_gnd_net_\,
            in3 => \N__11660\,
            lcout => \Lab_UT.scdp.b2a1.N_220_i\,
            ltout => \Lab_UT.scdp.b2a1.N_220_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.b2a1.asciiHex_2_i_o2_3_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111010"
        )
    port map (
            in0 => \N__10584\,
            in1 => \_gnd_net_\,
            in2 => \N__10563\,
            in3 => \N__12637\,
            lcout => \Lab_UT.scdp.N_282\,
            ltout => \Lab_UT.scdp.N_282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lsBitsi.q_esr_1_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__10555\,
            in1 => \_gnd_net_\,
            in2 => \N__10542\,
            in3 => \N__10538\,
            lcout => \Lab_UT.scdp.lsBitsD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21110\,
            ce => \N__11217\,
            sr => \N__20809\
        );

    \Lab_UT.scctrl.state_1_ret_5_RNI1UBG9_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001110"
        )
    port map (
            in0 => \N__11346\,
            in1 => \N__10526\,
            in2 => \N__20141\,
            in3 => \N__14000\,
            lcout => \Lab_UT.scctrl.sccLdLFSR\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lsBitsi.q_5_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10862\,
            in2 => \_gnd_net_\,
            in3 => \N__11231\,
            lcout => \Lab_UT.scdp.lsBitsi.lsBitsDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21101\,
            ce => 'H',
            sr => \N__20812\
        );

    \Lab_UT.scctrl.state_ret_13_RNI7RC32_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000100"
        )
    port map (
            in0 => \N__20114\,
            in1 => \N__10509\,
            in2 => \N__21723\,
            in3 => \N__23127\,
            lcout => \Lab_UT.scctrl.EmsLoaded\,
            ltout => \Lab_UT.scctrl.EmsLoaded_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNICOE1_0_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10503\,
            in3 => \N__21706\,
            lcout => \Lab_UT.sccElsBitsLd\,
            ltout => \Lab_UT.sccElsBitsLd_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lsBitsi.q_6_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10490\,
            in2 => \N__10500\,
            in3 => \N__10497\,
            lcout => \Lab_UT.scdp.lsBitsD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21101\,
            ce => 'H',
            sr => \N__20812\
        );

    \Lab_UT.scdp.lsBitsi.q_3_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__11232\,
            in1 => \N__10787\,
            in2 => \N__11697\,
            in3 => \N__10475\,
            lcout => \Lab_UT.scdp.lsBitsD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21101\,
            ce => 'H',
            sr => \N__20812\
        );

    \Lab_UT.scdp.msBitsi.q_esr_1_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010011000"
        )
    port map (
            in0 => \N__10630\,
            in1 => \N__10693\,
            in2 => \N__10724\,
            in3 => \N__11870\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21096\,
            ce => \N__11216\,
            sr => \N__20813\
        );

    \Lab_UT.scdp.msBitsi.q_esr_0_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010110100110"
        )
    port map (
            in0 => \N__11869\,
            in1 => \N__10715\,
            in2 => \N__10700\,
            in3 => \N__10629\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21096\,
            ce => \N__11216\,
            sr => \N__20813\
        );

    \Lab_UT.scdp.msBitsi.q_esr_2_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__10631\,
            in1 => \N__10694\,
            in2 => \N__10725\,
            in3 => \N__11871\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21096\,
            ce => \N__11216\,
            sr => \N__20813\
        );

    \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_1_1_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11059\,
            in1 => \N__12570\,
            in2 => \N__10743\,
            in3 => \N__11079\,
            lcout => \Lab_UT.scdp.b2a0.N_238_i\,
            ltout => \Lab_UT.scdp.b2a0.N_238_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_4_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010101011"
        )
    port map (
            in0 => \N__10696\,
            in1 => \N__10653\,
            in2 => \N__10728\,
            in3 => \N__11976\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21096\,
            ce => \N__11216\,
            sr => \N__20813\
        );

    \Lab_UT.scdp.msBitsi.q_esr_3_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10695\,
            in1 => \N__10722\,
            in2 => \_gnd_net_\,
            in3 => \N__10632\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21096\,
            ce => \N__11216\,
            sr => \N__20813\
        );

    \Lab_UT.scdp.msBitsi.q_esr_6_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001110"
        )
    port map (
            in0 => \N__10723\,
            in1 => \N__10652\,
            in2 => \N__10701\,
            in3 => \N__11975\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21096\,
            ce => \N__11216\,
            sr => \N__20813\
        );

    \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_0_1_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10651\,
            lcout => \Lab_UT.scdp.b2a0.N_224_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNI3LL8_0_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10617\,
            in1 => \N__10611\,
            in2 => \_gnd_net_\,
            in3 => \N__10828\,
            lcout => \Lab_UT.scdp.msBitsi.N_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8_1_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10829\,
            in1 => \N__10932\,
            in2 => \_gnd_net_\,
            in3 => \N__10926\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.msBitsi.N_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_1_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21709\,
            in2 => \N__10917\,
            in3 => \N__10974\,
            lcout => \ufifo.txdataDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21091\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNI7PL8_2_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10831\,
            in1 => \N__10902\,
            in2 => \_gnd_net_\,
            in3 => \N__10896\,
            lcout => \Lab_UT.scdp.msBitsi.N_1919_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNIBTL8_4_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10884\,
            in1 => \N__10878\,
            in2 => \_gnd_net_\,
            in3 => \N__10832\,
            lcout => \Lab_UT.scdp.msBitsi.N_1917_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNI2JO42_1_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__12088\,
            in1 => \N__12034\,
            in2 => \_gnd_net_\,
            in3 => \N__11971\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.N_332_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_5_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011101110"
        )
    port map (
            in0 => \N__10869\,
            in1 => \N__21710\,
            in2 => \N__10851\,
            in3 => \N__11552\,
            lcout => \ufifo.txdataDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21091\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNI019E_3_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__10830\,
            in1 => \_gnd_net_\,
            in2 => \N__10797\,
            in3 => \N__10788\,
            lcout => \Lab_UT.scdp.msBitsi.N_1915_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_3_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__10773\,
            in1 => \N__10764\,
            in2 => \N__21729\,
            in3 => \N__11085\,
            lcout => \ufifo.txdataDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_2_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__21707\,
            in1 => \N__11922\,
            in2 => \N__11022\,
            in3 => \N__11736\,
            lcout => \ufifo.txdataDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_4_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__10941\,
            in1 => \N__21708\,
            in2 => \N__10998\,
            in3 => \N__11094\,
            lcout => \ufifo.txdataDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNI4GMQ4_1_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110010110"
        )
    port map (
            in0 => \N__11846\,
            in1 => \N__11656\,
            in2 => \N__11628\,
            in3 => \N__11384\,
            lcout => \Lab_UT.scdp.N_552\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_esr_RNIA29D1_0_2_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12568\,
            in1 => \N__10965\,
            in2 => \N__11060\,
            in3 => \N__11074\,
            lcout => \Lab_UT.scdp.N_228_i_0\,
            ltout => \Lab_UT.scdp.N_228_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNI2TTL2_1_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__11623\,
            in1 => \N__11845\,
            in2 => \N__10968\,
            in3 => \N__11655\,
            lcout => \Lab_UT.scdp.u1.g0_0_i_a5_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_esr_RNIA29D1_2_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12569\,
            in1 => \N__10964\,
            in2 => \N__11061\,
            in3 => \N__11075\,
            lcout => \Lab_UT.scdp.N_228_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNI5V781_0_1_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12022\,
            in2 => \_gnd_net_\,
            in3 => \N__11955\,
            lcout => \Lab_UT.scdp.N_225_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNICF9Q4_7_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__11546\,
            in1 => \N__10953\,
            in2 => \N__11109\,
            in3 => \N__11792\,
            lcout => \Lab_UT.scdp.g0_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIPUDN_17_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11142\,
            in2 => \_gnd_net_\,
            in3 => \N__11034\,
            lcout => \Lab_UT.scdp.d2eData_3_0_1\,
            ltout => \Lab_UT.scdp.d2eData_3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNI116R2_1_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__11575\,
            in1 => \N__11621\,
            in2 => \N__10935\,
            in3 => \N__11840\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.u1.g0_0_i_a5_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNI7PSB8_0_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12717\,
            in1 => \N__11108\,
            in2 => \N__11097\,
            in3 => \N__11547\,
            lcout => \Lab_UT.scdp.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNIOKSG2_1_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__11841\,
            in1 => \N__11791\,
            in2 => \N__11661\,
            in3 => \N__11622\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.u1.g0_0_i_a5_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNIUCJ18_0_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12600\,
            in1 => \N__11459\,
            in2 => \N__11088\,
            in3 => \N__11548\,
            lcout => \Lab_UT.scdp.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIHOFN_22_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11136\,
            in2 => \_gnd_net_\,
            in3 => \N__11028\,
            lcout => \Lab_UT.scdp.d2eData_3_0_a2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNICL1I3_1_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110110111"
        )
    port map (
            in0 => \N__11963\,
            in1 => \N__12089\,
            in2 => \N__12048\,
            in3 => \N__11545\,
            lcout => \Lab_UT.scdp.N_276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_1_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17526\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21077\,
            ce => \N__12788\,
            sr => \N__20850\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_14_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13926\,
            lcout => \Lab_UT.scdp.prng_lfsr_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21077\,
            ce => \N__12788\,
            sr => \N__20850\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_17_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16890\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21077\,
            ce => \N__12788\,
            sr => \N__20850\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_22_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14103\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21077\,
            ce => \N__12788\,
            sr => \N__20850\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_25_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16851\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21077\,
            ce => \N__12788\,
            sr => \N__20850\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_3_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11415\,
            lcout => \Lab_UT.scdp.prng_lfsr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21077\,
            ce => \N__12788\,
            sr => \N__20850\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_30_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12501\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21077\,
            ce => \N__12788\,
            sr => \N__20850\
        );

    \Lab_UT.scctrl.state_1_RNO_9_0_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13223\,
            in2 => \_gnd_net_\,
            in3 => \N__22058\,
            lcout => \Lab_UT.scctrl.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.val_0_a2_3_3_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13541\,
            in1 => \N__17162\,
            in2 => \_gnd_net_\,
            in3 => \N__13031\,
            lcout => \Lab_UT.N_540i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.shifter_ret_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__11253\,
            in1 => \N__14526\,
            in2 => \_gnd_net_\,
            in3 => \N__15116\,
            lcout => \resetGen.N_243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21128\,
            ce => \N__13448\,
            sr => \N__20848\
        );

    \buart.Z_rx.shifter_ret_2_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18780\,
            lcout => \buart.bu_rx_data_i_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21123\,
            ce => \N__13446\,
            sr => \N__20842\
        );

    \Lab_UT.scctrl.shifter_ret_6_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18781\,
            in2 => \_gnd_net_\,
            in3 => \N__15084\,
            lcout => \Lab_UT.scctrl.N_534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21123\,
            ce => \N__13446\,
            sr => \N__20842\
        );

    \buart.Z_rx.shifter_1_5_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14900\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21123\,
            ce => \N__13446\,
            sr => \N__20842\
        );

    \buart.Z_rx.shifter_2_6_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14527\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21123\,
            ce => \N__13446\,
            sr => \N__20842\
        );

    \Lab_UT.scctrl.next_state_1_i_i_o2_5_0_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__13501\,
            in1 => \N__17161\,
            in2 => \_gnd_net_\,
            in3 => \N__15075\,
            lcout => \Lab_UT.scctrl.N_259i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_6_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11193\,
            in1 => \N__21721\,
            in2 => \_gnd_net_\,
            in3 => \N__11514\,
            lcout => \ufifo.txdataDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_5_RNIOMGF_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__18755\,
            in1 => \N__11172\,
            in2 => \_gnd_net_\,
            in3 => \N__12171\,
            lcout => \Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0\,
            ltout => \Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_1_RNI4BLT2_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18275\,
            in1 => \N__14522\,
            in2 => \N__11166\,
            in3 => \N__14380\,
            lcout => \Lab_UT.scctrl.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_9_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__22043\,
            in1 => \N__19731\,
            in2 => \N__22441\,
            in3 => \N__22292\,
            lcout => \Lab_UT.scctrl.N_415_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_8_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__22820\,
            in1 => \N__18065\,
            in2 => \N__15430\,
            in3 => \N__14632\,
            lcout => \Lab_UT.scctrl.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_4_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001010000"
        )
    port map (
            in0 => \N__11163\,
            in1 => \N__23202\,
            in2 => \N__11157\,
            in3 => \N__22970\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g1_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_1_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__12129\,
            in1 => \N__23690\,
            in2 => \N__11148\,
            in3 => \N__23507\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001010101010"
        )
    port map (
            in0 => \N__22542\,
            in1 => \N__14742\,
            in2 => \N__11145\,
            in3 => \N__15398\,
            lcout => \Lab_UT.scctrl.N_351_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txDataValidD_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13614\,
            in1 => \N__11493\,
            in2 => \_gnd_net_\,
            in3 => \N__13626\,
            lcout => \ufifo.txDataValidDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.un3_reset_count_i_o2_3_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__11249\,
            in1 => \N__14468\,
            in2 => \_gnd_net_\,
            in3 => \N__15079\,
            lcout => \N_243_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_0_RNIQM5P_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12974\,
            in1 => \N__13144\,
            in2 => \_gnd_net_\,
            in3 => \N__13170\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g1_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_0_RNIK3S32_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001000000"
        )
    port map (
            in0 => \N__15104\,
            in1 => \N__17827\,
            in2 => \N__11235\,
            in3 => \N__15180\,
            lcout => \Lab_UT.scctrl.g1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_fast_1_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart__rx_shifter_0_fast_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21102\,
            ce => \N__13441\,
            sr => \N__20830\
        );

    \buart.Z_rx.shifter_0_1_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12976\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21102\,
            ce => \N__13441\,
            sr => \N__20830\
        );

    \Lab_UT.scctrl.shifter_ret_0_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__13508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17155\,
            lcout => \Lab_UT.scctrl.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21102\,
            ce => \N__13441\,
            sr => \N__20830\
        );

    \buart.Z_rx.shifter_0_2_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13509\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21102\,
            ce => \N__13441\,
            sr => \N__20830\
        );

    \Lab_UT.scdp.msBitsi.q_esr_ctle_6_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16447\,
            in2 => \_gnd_net_\,
            in3 => \N__11230\,
            lcout => \Lab_UT.scdp.sccElsBitsLd_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_0_RNIDPMQ_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17128\,
            in1 => \N__12983\,
            in2 => \_gnd_net_\,
            in3 => \N__13171\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_0_RNI76D52_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000100000"
        )
    port map (
            in0 => \N__17855\,
            in1 => \N__15183\,
            in2 => \N__11394\,
            in3 => \N__15124\,
            lcout => \Lab_UT.scctrl.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_1_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22548\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_0_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__21724\,
            in1 => \N__11391\,
            in2 => \N__11373\,
            in3 => \N__12735\,
            lcout => \ufifo.txdataDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_5_RNIDAO06_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__23126\,
            in1 => \N__18278\,
            in2 => \N__20328\,
            in3 => \N__13984\,
            lcout => \Lab_UT.scctrl.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNIJOOS_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__20664\,
            in1 => \N__20118\,
            in2 => \_gnd_net_\,
            in3 => \N__21408\,
            lcout => \Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0dup_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIPVCP_4_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__13668\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13724\,
            lcout => \buart.Z_rx.sample_i_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.rddataDV.q_0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__13725\,
            in1 => \N__13669\,
            in2 => \N__11325\,
            in3 => \N__13860\,
            lcout => \Lab_UT.scdp.binVal_ValidD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21092\,
            ce => 'H',
            sr => \N__20816\
        );

    \buart.Z_rx.bitcount_es_RNIPVCP_2_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__13792\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13821\,
            lcout => \buart.Z_rx.N_230\,
            ltout => \buart.Z_rx.N_230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__13723\,
            in1 => \N__13667\,
            in2 => \N__11439\,
            in3 => \N__13859\,
            lcout => \N_232\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.k0h.q_2_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18574\,
            in1 => \N__16799\,
            in2 => \N__12587\,
            in3 => \N__12478\,
            lcout => \Lab_UT.scdp.key0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21092\,
            ce => 'H',
            sr => \N__20816\
        );

    \Lab_UT.scdp.k0h.q_3_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__12479\,
            in1 => \N__18576\,
            in2 => \N__11432\,
            in3 => \N__18533\,
            lcout => \Lab_UT.scdp.key0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21092\,
            ce => 'H',
            sr => \N__20816\
        );

    \Lab_UT.scdp.k0l.q_2_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18575\,
            in1 => \N__16800\,
            in2 => \N__11762\,
            in3 => \N__17555\,
            lcout => \Lab_UT.scdp.key0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21092\,
            ce => 'H',
            sr => \N__20816\
        );

    \Lab_UT.scdp.k0l.q_3_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__17556\,
            in1 => \N__18534\,
            in2 => \N__18623\,
            in3 => \N__11408\,
            lcout => \Lab_UT.scdp.key0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21092\,
            ce => 'H',
            sr => \N__20816\
        );

    \Lab_UT.scdp.rxdataD.q_1_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001001"
        )
    port map (
            in0 => \N__17051\,
            in1 => \N__17166\,
            in2 => \N__16641\,
            in3 => \N__13020\,
            lcout => \Lab_UT.scdp.binValD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21086\,
            ce => 'H',
            sr => \N__20819\
        );

    \Lab_UT.scdp.rxdataD.q_2_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__17165\,
            in1 => \N__13018\,
            in2 => \N__16639\,
            in3 => \N__17052\,
            lcout => \Lab_UT.scdp.binValD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21086\,
            ce => 'H',
            sr => \N__20819\
        );

    \Lab_UT.scdp.a2b.val_0_2_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__17050\,
            in1 => \N__17164\,
            in2 => \N__16640\,
            in3 => \N__13019\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.binVal_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_2_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__21593\,
            in1 => \N__12665\,
            in2 => \N__11397\,
            in3 => \N__21624\,
            lcout => \Lab_UT.scdp.u1.byteToDecryptZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21086\,
            ce => 'H',
            sr => \N__20819\
        );

    \Lab_UT.scdp.u1.q_1_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__21623\,
            in1 => \N__11502\,
            in2 => \N__21594\,
            in3 => \N__11617\,
            lcout => \Lab_UT.scdp.u1.byteToDecrypt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21086\,
            ce => 'H',
            sr => \N__20819\
        );

    \Lab_UT.scdp.a2b.val_i_1_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010010"
        )
    port map (
            in0 => \N__17163\,
            in1 => \N__13017\,
            in2 => \N__16638\,
            in3 => \N__17049\,
            lcout => \Lab_UT.scdp.N_73\,
            ltout => \Lab_UT.scdp.N_73_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_1_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12035\,
            in2 => \N__11496\,
            in3 => \N__16956\,
            lcout => \Lab_UT.scdp.byteToDecrypt_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21086\,
            ce => 'H',
            sr => \N__20819\
        );

    \Lab_UT.scctrl.r5.q_0_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21589\,
            in2 => \_gnd_net_\,
            in3 => \N__21622\,
            lcout => \Lab_UT.scctrl.delayload\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21086\,
            ce => 'H',
            sr => \N__20819\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_29_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12525\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21080\,
            ce => \N__12790\,
            sr => \N__20847\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_5_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12455\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21080\,
            ce => \N__12790\,
            sr => \N__20847\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_13_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17481\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21080\,
            ce => \N__12790\,
            sr => \N__20847\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIRBV41_5_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11445\,
            in1 => \N__11484\,
            in2 => \N__11478\,
            in3 => \N__11469\,
            lcout => \Lab_UT.scdp.d2eData_3_5\,
            ltout => \Lab_UT.scdp.d2eData_3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNI5V781_1_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11463\,
            in3 => \N__12021\,
            lcout => \Lab_UT.scdp.N_225_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_21_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14040\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21080\,
            ce => \N__12790\,
            sr => \N__20847\
        );

    \Lab_UT.scdp.u1.q_RNIOKSG2_0_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000101000"
        )
    port map (
            in0 => \N__12698\,
            in1 => \N__11962\,
            in2 => \N__12043\,
            in3 => \N__17267\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.u1.g0_0_i_a5_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNI3IJ18_0_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11579\,
            in1 => \N__11796\,
            in2 => \N__11745\,
            in3 => \N__11742\,
            lcout => \Lab_UT.scdp.N_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIT2EN_19_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11892\,
            in2 => \_gnd_net_\,
            in3 => \N__11667\,
            lcout => \Lab_UT.scdp.d2eData_3_0_3\,
            ltout => \Lab_UT.scdp.d2eData_3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI96HI1_3_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12830\,
            in1 => \N__11726\,
            in2 => \N__11730\,
            in3 => \N__16665\,
            lcout => \Lab_UT.scdp.N_255_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.b2a1.asciiHex_2_i_x2_3_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11727\,
            in1 => \N__12831\,
            in2 => \N__11718\,
            in3 => \N__11703\,
            lcout => \Lab_UT.scdp.N_226_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_19_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17430\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21078\,
            ce => \N__12789\,
            sr => \N__20851\
        );

    \Lab_UT.scdp.u1.q_RNIBG9H2_1_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \N__11830\,
            in1 => \N__11651\,
            in2 => \N__11627\,
            in3 => \N__12728\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.u1.N_539_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNIKMQ34_1_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11586\,
            in3 => \N__11574\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.N_426_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNI47LGA_1_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__12090\,
            in1 => \N__11544\,
            in2 => \N__11517\,
            in3 => \N__11775\,
            lcout => \Lab_UT.scdp.q_RNI47LGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_27_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17931\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21078\,
            ce => \N__12789\,
            sr => \N__20851\
        );

    \Lab_UT.scdp.b2a0.asciiHex_2_0_a2_0_x2_0_0_0_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12807\,
            in1 => \N__11805\,
            in2 => \N__11886\,
            in3 => \N__12861\,
            lcout => \Lab_UT.scdp.b2a0.N_258_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIK3K3_1_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12798\,
            in2 => \_gnd_net_\,
            in3 => \N__11853\,
            lcout => \Lab_UT.scdp.d2eData_3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIMSEN_20_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12837\,
            in2 => \_gnd_net_\,
            in3 => \N__12543\,
            lcout => \Lab_UT.scdp.d2eData_3_0_a2_0_4\,
            ltout => \Lab_UT.scdp.d2eData_3_0_a2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI0Q781_4_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12806\,
            in1 => \N__12860\,
            in2 => \N__11799\,
            in3 => \N__17310\,
            lcout => \Lab_UT.scdp.N_246_i\,
            ltout => \Lab_UT.scdp.N_246_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNI9Q034_1_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__12036\,
            in1 => \N__11769\,
            in2 => \N__11778\,
            in3 => \N__11972\,
            lcout => \Lab_UT.scdp.u0.L4_tx_data_0_a2_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNI41HI1_2_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12666\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12616\,
            lcout => \Lab_UT.scdp.N_256_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_2_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11763\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21072\,
            ce => \N__12785\,
            sr => \N__20853\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_10_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14058\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21072\,
            ce => \N__12785\,
            sr => \N__20853\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIO7U41_2_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12885\,
            in1 => \N__12105\,
            in2 => \N__12816\,
            in3 => \N__12099\,
            lcout => \Lab_UT.scdp.d2eData_3_2\,
            ltout => \Lab_UT.scdp.d2eData_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNI1L1F2_2_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111111111"
        )
    port map (
            in0 => \N__12667\,
            in1 => \_gnd_net_\,
            in2 => \N__12093\,
            in3 => \N__12081\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.g0_0_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNIGMI45_1_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110001"
        )
    port map (
            in0 => \N__12047\,
            in1 => \N__11988\,
            in2 => \N__11979\,
            in3 => \N__11973\,
            lcout => \Lab_UT.scdp.g0_0_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_2_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000001000000"
        )
    port map (
            in0 => \N__19131\,
            in1 => \N__15457\,
            in2 => \N__11901\,
            in3 => \N__23209\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g1_1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_0_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__19493\,
            in1 => \N__23524\,
            in2 => \N__11910\,
            in3 => \N__12375\,
            lcout => \Lab_UT.scctrl.g1_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_6_0_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__16151\,
            in1 => \N__11907\,
            in2 => \N__14661\,
            in3 => \N__22968\,
            lcout => \Lab_UT.scctrl.N_399_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_o2_9_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111011"
        )
    port map (
            in0 => \N__12165\,
            in1 => \N__14510\,
            in2 => \N__12188\,
            in3 => \N__18779\,
            lcout => \Lab_UT.scctrl.N_266i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_5_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__12891\,
            in1 => \N__19728\,
            in2 => \N__14660\,
            in3 => \N__22967\,
            lcout => \Lab_UT.scctrl.g1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_10_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22966\,
            in1 => \N__18038\,
            in2 => \_gnd_net_\,
            in3 => \N__22041\,
            lcout => \Lab_UT.scctrl.N_319_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_5_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21370\,
            in1 => \N__14766\,
            in2 => \N__12141\,
            in3 => \N__22286\,
            lcout => \Lab_UT.scctrl.N_414_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNIVJ4S_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20585\,
            in2 => \_gnd_net_\,
            in3 => \N__21369\,
            lcout => \Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.state_1_ret_rep1_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rst_i_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_0_RNIJFLD2_0_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__22042\,
            in1 => \N__19725\,
            in2 => \N__22464\,
            in3 => \N__22285\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_415_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNII8KJ5_3_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__12117\,
            in1 => \N__23191\,
            in2 => \N__12120\,
            in3 => \N__22969\,
            lcout => \Lab_UT.scctrl.g1_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep2_RNITVAN_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__22791\,
            in1 => \N__14652\,
            in2 => \N__18086\,
            in3 => \N__15443\,
            lcout => \Lab_UT.scctrl.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNIIHUU_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__18905\,
            in1 => \N__22790\,
            in2 => \N__16316\,
            in3 => \N__18756\,
            lcout => \Lab_UT.scctrl.g0_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_2_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13030\,
            in2 => \_gnd_net_\,
            in3 => \N__18782\,
            lcout => \Lab_UT.scctrl.N_241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21106\,
            ce => \N__13447\,
            sr => \N__20844\
        );

    \Lab_UT.scctrl.shifter_ret_14_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12111\,
            in2 => \_gnd_net_\,
            in3 => \N__14520\,
            lcout => \Lab_UT.scctrl.N_263_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21106\,
            ce => \N__13447\,
            sr => \N__20844\
        );

    \buart.Z_rx.shifter_ret_1_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17212\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21106\,
            ce => \N__13447\,
            sr => \N__20844\
        );

    \Lab_UT.scctrl.shifter_ret_5_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111011011101"
        )
    port map (
            in0 => \N__18783\,
            in1 => \N__12164\,
            in2 => \N__12192\,
            in3 => \N__14521\,
            lcout => \Lab_UT.scctrl.N_266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21106\,
            ce => \N__13447\,
            sr => \N__20844\
        );

    \buart.Z_rx.shifter_ret_0_rep1_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15083\,
            lcout => bu_rx_data_i_2_3_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21106\,
            ce => \N__13447\,
            sr => \N__20844\
        );

    \buart.Z_rx.shifter_0_4_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18784\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21106\,
            ce => \N__13447\,
            sr => \N__20844\
        );

    \Lab_UT.scdp.a2b.shifter_ret_RNISON11_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13747\,
            in1 => \N__15181\,
            in2 => \N__12924\,
            in3 => \N__15071\,
            lcout => \Lab_UT.scdp.a2b.val_0_tz_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.val_i_o2_0_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15072\,
            in1 => \N__13748\,
            in2 => \N__13517\,
            in3 => \N__15182\,
            lcout => \Lab_UT.scdp.a2b.N_280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_2_3_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15074\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21099\,
            ce => \N__13444\,
            sr => \N__20839\
        );

    \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_a2_3_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__17129\,
            in1 => \N__13494\,
            in2 => \_gnd_net_\,
            in3 => \N__12150\,
            lcout => \Lab_UT.scctrl.N_472_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_4_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12984\,
            in2 => \_gnd_net_\,
            in3 => \N__18788\,
            lcout => \Lab_UT.scctrl.N_241_reti\,
            ltout => \Lab_UT.scctrl.N_241_reti_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_3_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12144\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scctrl.N_241_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21099\,
            ce => \N__13444\,
            sr => \N__20839\
        );

    \buart.Z_rx.shifter_ret_0_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15073\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21099\,
            ce => \N__13444\,
            sr => \N__20839\
        );

    \Lab_UT.scctrl.shifter_ret_12_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__14937\,
            in1 => \N__17743\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scctrl.N_233_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21094\,
            ce => \N__13443\,
            sr => \N__20832\
        );

    \Lab_UT.scctrl.shifter_ret_12_RNIE3JF_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__12216\,
            in1 => \N__13404\,
            in2 => \_gnd_net_\,
            in3 => \N__12207\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNI0FVE3_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__18904\,
            in1 => \N__12201\,
            in2 => \N__12195\,
            in3 => \N__14338\,
            lcout => \Lab_UT.scctrl.N_351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_8_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17748\,
            in3 => \N__14936\,
            lcout => \Lab_UT.N_252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21094\,
            ce => \N__13443\,
            sr => \N__20832\
        );

    \buart.Z_rx.shifter_ret_3_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14938\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21094\,
            ce => \N__13443\,
            sr => \N__20832\
        );

    \buart.Z_rx.shifter_1_7_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21094\,
            ce => \N__13443\,
            sr => \N__20832\
        );

    \buart.Z_rx.shifter_2_fast_6_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14470\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart__rx_shifter_2_fast_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21094\,
            ce => \N__13443\,
            sr => \N__20832\
        );

    \buart.Z_rx.shifter_ret_5_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14469\,
            lcout => bu_rx_data_i_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21094\,
            ce => \N__13443\,
            sr => \N__20832\
        );

    \buart.Z_rx.bitcount_es_1_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__17694\,
            in1 => \N__13888\,
            in2 => \N__12240\,
            in3 => \N__13677\,
            lcout => \buart__rx_bitcount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21089\,
            ce => \N__12429\,
            sr => \N__20840\
        );

    \buart.Z_rx.bitcount_es_2_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__13889\,
            in1 => \N__17697\,
            in2 => \N__12228\,
            in3 => \N__13794\,
            lcout => \buart.Z_rx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21089\,
            ce => \N__12429\,
            sr => \N__20840\
        );

    \CONSTANT_ONE_LUT4_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => \CONSTANT_ONE_NET_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__13887\,
            in1 => \N__17696\,
            in2 => \N__12360\,
            in3 => \N__13865\,
            lcout => \buart.Z_rx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21089\,
            ce => \N__12429\,
            sr => \N__20840\
        );

    \buart.Z_rx.bitcount_es_3_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__17695\,
            in1 => \N__13890\,
            in2 => \N__13827\,
            in3 => \N__12441\,
            lcout => \buart.Z_rx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21089\,
            ce => \N__12429\,
            sr => \N__20840\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIQ8IQ3_0_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12357\,
            in1 => \N__12345\,
            in2 => \_gnd_net_\,
            in3 => \N__12330\,
            lcout => utb_txdata_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13861\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13676\,
            in2 => \_gnd_net_\,
            in3 => \N__12231\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13793\,
            in2 => \_gnd_net_\,
            in3 => \N__12219\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13822\,
            in2 => \_gnd_net_\,
            in3 => \N__12435\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_4_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__13886\,
            in1 => \N__17675\,
            in2 => \N__13731\,
            in3 => \N__12432\,
            lcout => \buart__rx_bitcount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21083\,
            ce => \N__12425\,
            sr => \N__20843\
        );

    \Lab_UT.scctrl.shifter_ret_3_RNIRA8MC_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__12389\,
            in1 => \N__12399\,
            in2 => \N__15219\,
            in3 => \N__16736\,
            lcout => \Lab_UT.scctrl.next_state_rst_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_1_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__22187\,
            in1 => \N__22424\,
            in2 => \N__22059\,
            in3 => \N__22827\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_418_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI91NK6_0_2_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__16703\,
            in1 => \N__19151\,
            in2 => \N__12402\,
            in3 => \N__23197\,
            lcout => \Lab_UT.scctrl.g0_2\,
            ltout => \Lab_UT.scctrl.g0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_3_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__16737\,
            in1 => \N__15218\,
            in2 => \N__12393\,
            in3 => \N__12390\,
            lcout => \Lab_UT.scctrl.next_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21079\,
            ce => \N__20900\,
            sr => \N__20849\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_7_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100010"
        )
    port map (
            in0 => \N__22828\,
            in1 => \N__22050\,
            in2 => \N__22454\,
            in3 => \N__22186\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_418_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_3_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__22188\,
            in1 => \N__14292\,
            in2 => \N__12378\,
            in3 => \N__21514\,
            lcout => \Lab_UT.scctrl.g1_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI6V451_2_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__22829\,
            in1 => \N__19152\,
            in2 => \N__21417\,
            in3 => \N__22051\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_39_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI6EDGH_2_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__12480\,
            in1 => \_gnd_net_\,
            in2 => \N__12363\,
            in3 => \N__15504\,
            lcout => \Lab_UT.state_1_RNI6EDGH_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_7_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17043\,
            in1 => \N__17885\,
            in2 => \N__18395\,
            in3 => \N__16157\,
            lcout => \Lab_UT.scctrl.N_404_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNI9TOB1_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__18356\,
            in1 => \N__20657\,
            in2 => \_gnd_net_\,
            in3 => \N__22052\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_22_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNI9C1NH_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15503\,
            in2 => \N__12531\,
            in3 => \N__12511\,
            lcout => \Lab_UT.state_1_ret_0_RNI9C1NH_0\,
            ltout => \Lab_UT.state_1_ret_0_RNI9C1NH_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.k3h.q_0_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__17617\,
            in1 => \N__12848\,
            in2 => \N__12528\,
            in3 => \N__18664\,
            lcout => \Lab_UT.scdp.key3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21076\,
            ce => 'H',
            sr => \N__20820\
        );

    \Lab_UT.scdp.k3h.q_1_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__17374\,
            in1 => \N__12524\,
            in2 => \N__18689\,
            in3 => \N__12512\,
            lcout => \Lab_UT.scdp.key3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21076\,
            ce => 'H',
            sr => \N__20820\
        );

    \Lab_UT.scdp.k3h.q_2_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__12513\,
            in1 => \N__18660\,
            in2 => \N__12497\,
            in3 => \N__16801\,
            lcout => \Lab_UT.scdp.key3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21076\,
            ce => 'H',
            sr => \N__20820\
        );

    \Lab_UT.scdp.k0h.q_0_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18658\,
            in1 => \N__17616\,
            in2 => \N__12878\,
            in3 => \N__12476\,
            lcout => \Lab_UT.scdp.key0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21076\,
            ce => 'H',
            sr => \N__20820\
        );

    \Lab_UT.scdp.k0h.q_1_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__12477\,
            in1 => \N__18659\,
            in2 => \N__12456\,
            in3 => \N__17375\,
            lcout => \Lab_UT.scdp.key0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21076\,
            ce => 'H',
            sr => \N__20820\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_24_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16869\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21074\,
            ce => \N__12787\,
            sr => \N__20852\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_0_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17577\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21074\,
            ce => \N__12787\,
            sr => \N__20852\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_16_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16908\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21074\,
            ce => \N__12787\,
            sr => \N__20852\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI9U1R_0_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12759\,
            in1 => \N__12537\,
            in2 => \N__12753\,
            in3 => \N__12744\,
            lcout => \Lab_UT.scdp.d2eData_3_0\,
            ltout => \Lab_UT.scdp.d2eData_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNIJLK81_0_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12738\,
            in3 => \N__17262\,
            lcout => \Lab_UT.scdp.N_262_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNINM5R2_0_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001100000"
        )
    port map (
            in0 => \N__12626\,
            in1 => \N__12671\,
            in2 => \N__17268\,
            in3 => \N__12691\,
            lcout => \Lab_UT.scdp.u1.g0_0_i_a5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNINM5R2_0_0_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001100000"
        )
    port map (
            in0 => \N__12690\,
            in1 => \N__17263\,
            in2 => \N__12672\,
            in3 => \N__12625\,
            lcout => \Lab_UT.scdp.u1.g0_0_i_a5_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_6_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12591\,
            lcout => \Lab_UT.scdp.prng_lfsr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21071\,
            ce => \N__12786\,
            sr => \N__20854\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_20_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14087\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21071\,
            ce => \N__12786\,
            sr => \N__20854\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_8_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14132\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21071\,
            ce => \N__12786\,
            sr => \N__20854\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_18_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14072\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21071\,
            ce => \N__12786\,
            sr => \N__20854\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_4_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12879\,
            lcout => \Lab_UT.scdp.prng_lfsr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21071\,
            ce => \N__12786\,
            sr => \N__20854\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_28_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12852\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21071\,
            ce => \N__12786\,
            sr => \N__20854\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_11_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14117\,
            lcout => \Lab_UT.scdp.prng_lfsr_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21071\,
            ce => \N__12786\,
            sr => \N__20854\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_26_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16776\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21071\,
            ce => \N__12786\,
            sr => \N__20854\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_12_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14018\,
            lcout => \Lab_UT.scdp.prng_lfsr_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21070\,
            ce => \N__12784\,
            sr => \N__20856\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_9_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17334\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21070\,
            ce => \N__12784\,
            sr => \N__20856\
        );

    \Lab_UT.scctrl.sccEldByte_i_a2_0_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12914\,
            in1 => \N__12897\,
            in2 => \N__13549\,
            in3 => \N__18803\,
            lcout => \Lab_UT.scctrl.N_385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_a2_2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18804\,
            in2 => \_gnd_net_\,
            in3 => \N__15106\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_534_reti_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_7_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13047\,
            in3 => \N__13044\,
            lcout => \Lab_UT.scctrl.N_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21137\,
            ce => \N__13449\,
            sr => \N__20855\
        );

    \Lab_UT.scdp.a2b.shifter_ret_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17213\,
            in2 => \N__13550\,
            in3 => \N__13037\,
            lcout => \Lab_UT.N_540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21137\,
            ce => \N__13449\,
            sr => \N__20855\
        );

    \Lab_UT.scctrl.shifter_ret_13_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011001110110011"
        )
    port map (
            in0 => \N__15107\,
            in1 => \N__13537\,
            in2 => \N__17217\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scctrl.N_259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21137\,
            ce => \N__13449\,
            sr => \N__20855\
        );

    \Lab_UT.scctrl.state_1_RNO_8_0_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__16158\,
            in1 => \N__14514\,
            in2 => \_gnd_net_\,
            in3 => \N__13411\,
            lcout => \Lab_UT.scctrl.g0_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_2_0_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__12903\,
            in1 => \N__18245\,
            in2 => \N__18441\,
            in3 => \N__15455\,
            lcout => \Lab_UT.scctrl.g0_1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.sccEldByte_i_a2_0_1_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14926\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15105\,
            lcout => \Lab_UT.scctrl.sccEldByte_i_a2_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_10_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20577\,
            in2 => \_gnd_net_\,
            in3 => \N__21314\,
            lcout => \Lab_UT.scctrl.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_9_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22034\,
            in1 => \N__18039\,
            in2 => \_gnd_net_\,
            in3 => \N__22975\,
            lcout => \Lab_UT.scctrl.N_319_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_1_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__13083\,
            in1 => \N__23706\,
            in2 => \N__23529\,
            in3 => \N__13065\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_1_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111111111"
        )
    port map (
            in0 => \N__13104\,
            in1 => \_gnd_net_\,
            in2 => \N__13098\,
            in3 => \N__15456\,
            lcout => \Lab_UT.scctrl.N_235_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_3_RNIUPHA1_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16576\,
            in1 => \N__13258\,
            in2 => \N__14939\,
            in3 => \N__14850\,
            lcout => \Lab_UT.scctrl.N_444_0\,
            ltout => \Lab_UT.scctrl.N_444_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_8_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110010"
        )
    port map (
            in0 => \N__13355\,
            in1 => \N__15197\,
            in2 => \N__13095\,
            in3 => \N__15069\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_223_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_4_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22268\,
            in1 => \N__13092\,
            in2 => \N__13086\,
            in3 => \N__21316\,
            lcout => \Lab_UT.scctrl.N_414_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.state_1_ret_fast_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22580\,
            lcout => rst_i_fast,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNO_4_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111101100"
        )
    port map (
            in0 => \N__15070\,
            in1 => \N__13077\,
            in2 => \N__15201\,
            in3 => \N__13356\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_223_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNO_3_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21317\,
            in1 => \N__18099\,
            in2 => \N__13071\,
            in3 => \N__22269\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_414_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNO_1_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__23696\,
            in1 => \N__23525\,
            in2 => \N__13068\,
            in3 => \N__13061\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__15447\,
            in1 => \_gnd_net_\,
            in2 => \N__13050\,
            in3 => \N__15804\,
            lcout => \Lab_UT.scctrl.N_235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep1_RNIEMAA2_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__16149\,
            in1 => \N__13116\,
            in2 => \N__20529\,
            in3 => \N__13128\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep1_RNIKQNN6_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__23149\,
            in1 => \N__13953\,
            in2 => \N__13122\,
            in3 => \N__19316\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_0_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep2_RNI4KGMF_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001111"
        )
    port map (
            in0 => \N__14653\,
            in1 => \N__14232\,
            in2 => \N__13119\,
            in3 => \N__19376\,
            lcout => \Lab_UT.scctrl.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNO_5_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001000"
        )
    port map (
            in0 => \N__20528\,
            in1 => \N__16150\,
            in2 => \N__13200\,
            in3 => \N__22944\,
            lcout => \Lab_UT.scctrl.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_2_RNI2SHF_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13399\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16148\,
            lcout => \Lab_UT.scctrl.N_487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_2_RNI8G3S_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__13250\,
            in1 => \N__13398\,
            in2 => \_gnd_net_\,
            in3 => \N__16988\,
            lcout => \Lab_UT.scctrl.N_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_15_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__16989\,
            in1 => \N__16147\,
            in2 => \N__13259\,
            in3 => \N__15878\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_2_0_0_a3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_13_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15952\,
            in1 => \N__14482\,
            in2 => \N__13110\,
            in3 => \N__14371\,
            lcout => \Lab_UT.scctrl.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_13_RNIORKJ_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13219\,
            in2 => \_gnd_net_\,
            in3 => \N__21873\,
            lcout => \Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0\,
            ltout => \Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep1_RNI5JDF1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__20521\,
            in1 => \N__19603\,
            in2 => \N__13107\,
            in3 => \N__16099\,
            lcout => \Lab_UT.scctrl.N_399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_2_RNI1JJ81_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__16990\,
            in1 => \N__13254\,
            in2 => \N__19608\,
            in3 => \N__13400\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_i_o7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep2_RNIE3HB2_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__14592\,
            in1 => \N__13272\,
            in2 => \N__13266\,
            in3 => \N__16100\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_12_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep2_RNIBDOL6_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__13185\,
            in1 => \N__14208\,
            in2 => \N__13263\,
            in3 => \N__23128\,
            lcout => \Lab_UT.scctrl.g0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNO_6_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__21875\,
            in1 => \N__13260\,
            in2 => \N__13224\,
            in3 => \N__16991\,
            lcout => \Lab_UT.scctrl.g0_1_i_a8_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNIBUL06_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21391\,
            in1 => \N__22250\,
            in2 => \N__20661\,
            in3 => \N__21479\,
            lcout => \Lab_UT.scctrl.N_401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNIQILS_0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__21874\,
            in1 => \N__19890\,
            in2 => \_gnd_net_\,
            in3 => \N__18265\,
            lcout => \Lab_UT.scctrl.N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_9_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__15092\,
            in1 => \N__13179\,
            in2 => \_gnd_net_\,
            in3 => \N__15169\,
            lcout => \Lab_UT.scctrl.N_12_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_11_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13173\,
            in1 => \N__13148\,
            in2 => \_gnd_net_\,
            in3 => \N__13563\,
            lcout => \Lab_UT.scctrl.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_0_RNI51T61_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__13313\,
            in1 => \N__13172\,
            in2 => \N__13149\,
            in3 => \N__13562\,
            lcout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0\,
            ltout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110011000"
        )
    port map (
            in0 => \N__15168\,
            in1 => \N__15091\,
            in2 => \N__13359\,
            in3 => \N__13324\,
            lcout => \Lab_UT.scctrl.N_223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_1_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010101110"
        )
    port map (
            in0 => \N__13325\,
            in1 => \N__13345\,
            in2 => \N__15120\,
            in3 => \N__15170\,
            lcout => \Lab_UT.scctrl.N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110011000"
        )
    port map (
            in0 => \N__15171\,
            in1 => \N__15096\,
            in2 => \N__13354\,
            in3 => \N__13326\,
            lcout => \Lab_UT.scctrl.N_223_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_3_RNIESH11_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16241\,
            in1 => \N__14836\,
            in2 => \N__13314\,
            in3 => \N__13332\,
            lcout => \Lab_UT.scctrl.N_444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_ret_0_fast_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15097\,
            lcout => bu_rx_data_i_2_fast_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21103\,
            ce => \N__13445\,
            sr => \N__20836\
        );

    \Lab_UT.scctrl.shifter_ret_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13290\,
            in2 => \_gnd_net_\,
            in3 => \N__13302\,
            lcout => \Lab_UT.scctrl.N_271_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21098\,
            ce => \N__13442\,
            sr => \N__20845\
        );

    \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_5_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13545\,
            in2 => \_gnd_net_\,
            in3 => \N__17196\,
            lcout => \Lab_UT.scctrl.N_219i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_RNI4H6R_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__13716\,
            in1 => \N__13670\,
            in2 => \N__13284\,
            in3 => \N__13412\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_RNI7U912_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13275\,
            in3 => \N__13764\,
            lcout => \N_272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_fast_0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17197\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart__rx_shifter_1_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21098\,
            ce => \N__13442\,
            sr => \N__20845\
        );

    \buart.Z_rx.shifter_0_fast_2_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13547\,
            lcout => \buart__rx_shifter_0_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21098\,
            ce => \N__13442\,
            sr => \N__20845\
        );

    \buart.Z_rx.shifter_ret_4_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__13546\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21098\,
            ce => \N__13442\,
            sr => \N__20845\
        );

    \buart.Z_rx.shifter_1_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17198\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21098\,
            ce => \N__13442\,
            sr => \N__20845\
        );

    \Lab_UT.scctrl.sccEldByte_i_o2_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__13673\,
            in1 => \N__14475\,
            in2 => \N__13730\,
            in3 => \N__13766\,
            lcout => \Lab_UT.scctrl.N_284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIPVCP_0_2_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__13791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13820\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcountN11_15_i_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_0_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__13858\,
            in1 => \N__13726\,
            in2 => \N__13416\,
            in3 => \N__13675\,
            lcout => \buart.Z_rx.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_2_RNI4KBA1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__14474\,
            in1 => \N__13672\,
            in2 => \N__16146\,
            in3 => \N__13413\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_70_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13721\,
            in1 => \N__13765\,
            in2 => \N__13362\,
            in3 => \N__15902\,
            lcout => \Lab_UT.scctrl.next_state_rst_0_3_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIOP0V3_4_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001111"
        )
    port map (
            in0 => \N__13767\,
            in1 => \N__13722\,
            in2 => \N__17791\,
            in3 => \N__13674\,
            lcout => \buart.Z_rx.N_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNI3D361_2_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__13857\,
            in1 => \_gnd_net_\,
            in2 => \N__13826\,
            in3 => \N__13790\,
            lcout => \buart__rx_N_86_i_0_o2_1_0\,
            ltout => \buart__rx_N_86_i_0_o2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_8_RNIG4702_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__13749\,
            in1 => \N__13717\,
            in2 => \N__13680\,
            in3 => \N__13671\,
            lcout => \Lab_UT.scctrl.N_261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.r4.q_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13610\,
            lcout => \Lab_UT.scctrl.r4.delay4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21087\,
            ce => 'H',
            sr => \N__20821\
        );

    \Lab_UT.scctrl.r3.q_0_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13590\,
            lcout => \Lab_UT.scctrl.delay3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21087\,
            ce => 'H',
            sr => \N__20821\
        );

    \Lab_UT.scctrl.r1.q_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15920\,
            in1 => \N__13584\,
            in2 => \N__21728\,
            in3 => \N__13578\,
            lcout => \Lab_UT.scctrl.delay1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21087\,
            ce => 'H',
            sr => \N__20821\
        );

    \Lab_UT.scctrl.r2.q_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13596\,
            lcout => \Lab_UT.scctrl.delay2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21087\,
            ce => 'H',
            sr => \N__20821\
        );

    \Lab_UT.scctrl.sccEldByte_i_a2_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16138\,
            in2 => \_gnd_net_\,
            in3 => \N__15196\,
            lcout => \Lab_UT.scctrl.N_384\,
            ltout => \Lab_UT.scctrl.N_384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNIRGEB5_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13577\,
            in1 => \N__15919\,
            in2 => \N__13566\,
            in3 => \N__21717\,
            lcout => OPEN,
            ltout => \Lab_UT.N_100_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u2.q_esr_ctle_7_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13908\,
            in3 => \N__20862\,
            lcout => \Lab_UT.scdp.u2.N_100_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_15_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14633\,
            in1 => \N__17036\,
            in2 => \N__17896\,
            in3 => \N__16152\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_8_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13896\,
            in3 => \N__19331\,
            lcout => \Lab_UT.scctrl.G_24_i_o7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_5_0_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14634\,
            in1 => \N__17037\,
            in2 => \N__17894\,
            in3 => \N__16153\,
            lcout => \Lab_UT.scctrl.N_404_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_7_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100010"
        )
    port map (
            in0 => \N__22819\,
            in1 => \N__22054\,
            in2 => \N__22462\,
            in3 => \N__22209\,
            lcout => \Lab_UT.scctrl.N_418_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNO_4_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14636\,
            in1 => \N__17042\,
            in2 => \N__17895\,
            in3 => \N__16156\,
            lcout => \Lab_UT.scctrl.N_404_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_5_RNO_3_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16154\,
            in1 => \N__17884\,
            in2 => \N__17053\,
            in3 => \N__14635\,
            lcout => \Lab_UT.scctrl.N_404_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNO_4_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14637\,
            in1 => \N__17041\,
            in2 => \N__17897\,
            in3 => \N__16155\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_404_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNO_1_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__13944\,
            in1 => \N__19332\,
            in2 => \N__13893\,
            in3 => \N__21497\,
            lcout => \Lab_UT.scctrl.g0_2_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_3_RNI216C3_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15460\,
            in2 => \_gnd_net_\,
            in3 => \N__21495\,
            lcout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0\,
            ltout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_0_RNIIKTO3_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__22046\,
            in1 => \_gnd_net_\,
            in2 => \N__14004\,
            in3 => \N__19729\,
            lcout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNI71T5A_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__15534\,
            in1 => \N__22199\,
            in2 => \N__14001\,
            in3 => \N__13968\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI0F8BG_0_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__22201\,
            in1 => \N__21411\,
            in2 => \N__13962\,
            in3 => \N__13959\,
            lcout => \Lab_UT.scctrl.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNIQILS_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22045\,
            in2 => \N__19906\,
            in3 => \N__18264\,
            lcout => \Lab_UT.scctrl.N_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNO_3_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__22200\,
            in1 => \N__20655\,
            in2 => \_gnd_net_\,
            in3 => \N__21410\,
            lcout => \Lab_UT.scctrl.g0_8_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNO_3_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__21412\,
            in1 => \N__20656\,
            in2 => \_gnd_net_\,
            in3 => \N__22202\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNO_1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__21496\,
            in1 => \N__13938\,
            in2 => \N__13929\,
            in3 => \N__19333\,
            lcout => \Lab_UT.scctrl.g0_2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.k1h.q_2_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18665\,
            in1 => \N__16820\,
            in2 => \N__13925\,
            in3 => \N__17505\,
            lcout => \Lab_UT.scdp.key1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21075\,
            ce => 'H',
            sr => \N__20824\
        );

    \Lab_UT.scdp.k1h.q_3_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__17506\,
            in1 => \N__18668\,
            in2 => \N__14150\,
            in3 => \N__18531\,
            lcout => \Lab_UT.scdp.key1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21075\,
            ce => 'H',
            sr => \N__20824\
        );

    \Lab_UT.scdp.k1l.q_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18666\,
            in1 => \N__17626\,
            in2 => \N__14133\,
            in3 => \N__17354\,
            lcout => \Lab_UT.scdp.key1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21075\,
            ce => 'H',
            sr => \N__20824\
        );

    \Lab_UT.scdp.k1l.q_3_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__17356\,
            in1 => \N__18669\,
            in2 => \N__14118\,
            in3 => \N__18532\,
            lcout => \Lab_UT.scdp.key1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21075\,
            ce => 'H',
            sr => \N__20824\
        );

    \Lab_UT.scdp.k2h.q_2_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__18483\,
            in1 => \N__14099\,
            in2 => \N__18690\,
            in3 => \N__16824\,
            lcout => \Lab_UT.scdp.key2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21075\,
            ce => 'H',
            sr => \N__20824\
        );

    \Lab_UT.scdp.k2h.q_0_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17627\,
            in1 => \N__18670\,
            in2 => \N__14088\,
            in3 => \N__18482\,
            lcout => \Lab_UT.scdp.key2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21075\,
            ce => 'H',
            sr => \N__20824\
        );

    \Lab_UT.scdp.k2l.q_2_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18667\,
            in1 => \N__16825\,
            in2 => \N__14073\,
            in3 => \N__17455\,
            lcout => \Lab_UT.scdp.key2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21075\,
            ce => 'H',
            sr => \N__20824\
        );

    \Lab_UT.scdp.k1l.q_2_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__17355\,
            in1 => \N__14051\,
            in2 => \N__16827\,
            in3 => \N__18674\,
            lcout => \Lab_UT.scdp.key1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21075\,
            ce => 'H',
            sr => \N__20824\
        );

    \Lab_UT.scdp.k2h.q_1_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__18489\,
            in1 => \N__18688\,
            in2 => \N__14036\,
            in3 => \N__17402\,
            lcout => \Lab_UT.scdp.key2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21073\,
            ce => 'H',
            sr => \N__20827\
        );

    \Lab_UT.scdp.k1h.q_0_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18687\,
            in1 => \N__17628\,
            in2 => \N__14019\,
            in3 => \N__17507\,
            lcout => \Lab_UT.scdp.key1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21073\,
            ce => 'H',
            sr => \N__20827\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_16_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20354\,
            in1 => \N__15747\,
            in2 => \_gnd_net_\,
            in3 => \N__16280\,
            lcout => \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_8_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__14631\,
            in1 => \N__23453\,
            in2 => \N__18071\,
            in3 => \N__22804\,
            lcout => \Lab_UT.scctrl.N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_3_0_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010000"
        )
    port map (
            in0 => \N__18263\,
            in1 => \N__19392\,
            in2 => \N__14196\,
            in3 => \N__23190\,
            lcout => \Lab_UT.scctrl.g0_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep2_RNIN4FF_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__14630\,
            in1 => \N__18004\,
            in2 => \_gnd_net_\,
            in3 => \N__22803\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g1_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIVOU53_3_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010100000"
        )
    port map (
            in0 => \N__15461\,
            in1 => \N__23189\,
            in2 => \N__14175\,
            in3 => \N__22971\,
            lcout => \Lab_UT.scctrl.g1_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_14_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__21305\,
            in1 => \N__16305\,
            in2 => \N__20605\,
            in3 => \N__14172\,
            lcout => \Lab_UT.scctrl.next_state_rst_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_0_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14516\,
            in1 => \N__15896\,
            in2 => \N__15977\,
            in3 => \N__14384\,
            lcout => \Lab_UT.scctrl.N_290\,
            ltout => \Lab_UT.scctrl.N_290_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNO_2_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__18437\,
            in1 => \_gnd_net_\,
            in2 => \N__14166\,
            in3 => \N__18238\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNO_0_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__20284\,
            in1 => \N__23496\,
            in2 => \N__14163\,
            in3 => \N__14259\,
            lcout => \Lab_UT.scctrl.next_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_4_0_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111111111"
        )
    port map (
            in0 => \N__14385\,
            in1 => \N__14160\,
            in2 => \N__15903\,
            in3 => \N__18438\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_0_0_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18702\,
            in1 => \N__14226\,
            in2 => \N__14220\,
            in3 => \N__14217\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_0_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__23497\,
            in1 => \N__20285\,
            in2 => \N__14211\,
            in3 => \N__20183\,
            lcout => \Lab_UT.scctrl.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21138\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_0_RNIJFLD2_1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__22031\,
            in1 => \N__19712\,
            in2 => \N__22420\,
            in3 => \N__22267\,
            lcout => \Lab_UT.scctrl.N_415_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNO_3_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001100110011"
        )
    port map (
            in0 => \N__18787\,
            in1 => \N__23572\,
            in2 => \N__18903\,
            in3 => \N__22700\,
            lcout => \Lab_UT.scctrl.g0_1_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNISO7C1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__22698\,
            in1 => \N__18887\,
            in2 => \N__23589\,
            in3 => \N__18785\,
            lcout => \Lab_UT.scctrl.g0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_7_0_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19847\,
            in2 => \_gnd_net_\,
            in3 => \N__22033\,
            lcout => \Lab_UT.scctrl.g3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep1_RNICQA1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__18203\,
            in1 => \N__20522\,
            in2 => \_gnd_net_\,
            in3 => \N__16306\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNIBVSV_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__18786\,
            in1 => \N__18897\,
            in2 => \N__14184\,
            in3 => \N__22699\,
            lcout => \Lab_UT.scctrl.next_state_rst_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNO_4_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011100"
        )
    port map (
            in0 => \N__22032\,
            in1 => \N__18231\,
            in2 => \N__19873\,
            in3 => \N__23187\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_1_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNO_1_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14181\,
            in1 => \N__14268\,
            in2 => \N__14262\,
            in3 => \N__19389\,
            lcout => \Lab_UT.scctrl.g0_1_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_12_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19315\,
            in2 => \_gnd_net_\,
            in3 => \N__14253\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_24_i_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_6_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__18406\,
            in1 => \N__19369\,
            in2 => \N__14244\,
            in3 => \N__14241\,
            lcout => \Lab_UT.scctrl.G_24_i_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_11_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20523\,
            in1 => \N__19577\,
            in2 => \_gnd_net_\,
            in3 => \N__19681\,
            lcout => \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNO_6_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14373\,
            in1 => \N__14518\,
            in2 => \N__15974\,
            in3 => \N__15892\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_290_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNO_2_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__18416\,
            in1 => \N__15695\,
            in2 => \N__14235\,
            in3 => \N__15543\,
            lcout => \Lab_UT.scctrl.g0_2_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNO_6_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14374\,
            in1 => \N__14519\,
            in2 => \N__15975\,
            in3 => \N__15891\,
            lcout => \Lab_UT.scctrl.N_290_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_1_RNI4BLT2_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14517\,
            in1 => \N__15879\,
            in2 => \N__18277\,
            in3 => \N__14372\,
            lcout => \Lab_UT.scctrl.N_8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI6O741_2_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__22741\,
            in1 => \N__15451\,
            in2 => \N__18433\,
            in3 => \N__19125\,
            lcout => \Lab_UT.scctrl.next_state_rst_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIECCO9_2_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__19132\,
            in1 => \N__14550\,
            in2 => \N__14541\,
            in3 => \N__23150\,
            lcout => \Lab_UT.scctrl.next_state_rst_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_5_RNI1VIJ5_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22284\,
            in1 => \N__16207\,
            in2 => \N__18058\,
            in3 => \N__21480\,
            lcout => \Lab_UT.scctrl.N_419_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep1_RNIHGED_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__19573\,
            in1 => \N__20508\,
            in2 => \_gnd_net_\,
            in3 => \N__19687\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNIDO8N1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__20643\,
            in1 => \N__23600\,
            in2 => \N__14544\,
            in3 => \N__21333\,
            lcout => \Lab_UT.scctrl.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_5_RNO_5_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15901\,
            in1 => \N__14515\,
            in2 => \N__15976\,
            in3 => \N__14370\,
            lcout => \Lab_UT.scctrl.N_290_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNO_6_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18028\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16206\,
            lcout => \Lab_UT.scctrl.g0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_fast_RNIKKMF_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__19572\,
            in1 => \N__15743\,
            in2 => \_gnd_net_\,
            in3 => \N__20350\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNIGSGP1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__20642\,
            in1 => \N__23599\,
            in2 => \N__14280\,
            in3 => \N__21332\,
            lcout => \Lab_UT.scctrl.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__15663\,
            in1 => \N__14277\,
            in2 => \N__15624\,
            in3 => \N__20037\,
            lcout => \Lab_UT.N_245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21112\,
            ce => 'H',
            sr => \N__20817\
        );

    \Lab_UT.scctrl.state_ret_12_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111110101011"
        )
    port map (
            in0 => \N__20038\,
            in1 => \N__23390\,
            in2 => \N__20287\,
            in3 => \N__14571\,
            lcout => \Lab_UT.scctrl.N_240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21112\,
            ce => 'H',
            sr => \N__20817\
        );

    \Lab_UT.scctrl.state_ret_RNI3VN3G_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__15257\,
            in1 => \N__15312\,
            in2 => \N__18355\,
            in3 => \N__15287\,
            lcout => \Lab_UT.scctrl.next_state_rst\,
            ltout => \Lab_UT.scctrl.next_state_rst_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_fast_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__20268\,
            in1 => \_gnd_net_\,
            in2 => \N__14664\,
            in3 => \N__23392\,
            lcout => \Lab_UT.scctrl.state_i_1_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21112\,
            ce => 'H',
            sr => \N__20817\
        );

    \Lab_UT.scctrl.state_ret_rep1_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__23389\,
            in1 => \N__20269\,
            in2 => \_gnd_net_\,
            in3 => \N__16353\,
            lcout => \Lab_UT.scctrl.state_i_1_0_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21112\,
            ce => 'H',
            sr => \N__20817\
        );

    \Lab_UT.scctrl.state_ret_5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__20039\,
            in1 => \N__20276\,
            in2 => \N__16359\,
            in3 => \N__23391\,
            lcout => \Lab_UT.scctrl.N_240_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21112\,
            ce => 'H',
            sr => \N__20817\
        );

    \Lab_UT.scctrl.state_ret_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__23388\,
            in1 => \N__20267\,
            in2 => \_gnd_net_\,
            in3 => \N__16352\,
            lcout => \Lab_UT.scctrl.state_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21112\,
            ce => 'H',
            sr => \N__20817\
        );

    \Lab_UT.scctrl.state_ret_rep2_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010100001111"
        )
    port map (
            in0 => \N__16354\,
            in1 => \_gnd_net_\,
            in2 => \N__20286\,
            in3 => \N__23393\,
            lcout => \Lab_UT.scctrl.state_i_1_0_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21112\,
            ce => 'H',
            sr => \N__20817\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001110101100"
        )
    port map (
            in0 => \N__14805\,
            in1 => \N__19496\,
            in2 => \N__23452\,
            in3 => \N__20015\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_299_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__20184\,
            in1 => \N__15620\,
            in2 => \N__14574\,
            in3 => \N__14556\,
            lcout => \Lab_UT_scctrl_N_223_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21104\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNI09OAV_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001101"
        )
    port map (
            in0 => \N__23352\,
            in1 => \N__14570\,
            in2 => \N__20283\,
            in3 => \N__20014\,
            lcout => \Lab_UT.scctrl.N_240_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_7_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__15792\,
            in1 => \N__15702\,
            in2 => \_gnd_net_\,
            in3 => \N__23351\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_2_0_0_a3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_3_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22842\,
            in1 => \N__14796\,
            in2 => \N__14715\,
            in3 => \N__14712\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_24_i_a3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_1_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111111"
        )
    port map (
            in0 => \N__20016\,
            in1 => \N__14685\,
            in2 => \N__14703\,
            in3 => \N__14700\,
            lcout => \Lab_UT.scctrl.N_398i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__22841\,
            in1 => \N__14789\,
            in2 => \N__14694\,
            in3 => \N__22192\,
            lcout => \Lab_UT.scctrl.G_24_i_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_5_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__19495\,
            in1 => \N__20258\,
            in2 => \_gnd_net_\,
            in3 => \N__23350\,
            lcout => \Lab_UT.scctrl.G_24_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_4_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__16365\,
            in1 => \N__14778\,
            in2 => \N__19008\,
            in3 => \N__14790\,
            lcout => \Lab_UT.scctrl.N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI9JP5A_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101000"
        )
    port map (
            in0 => \N__22189\,
            in1 => \N__22027\,
            in2 => \N__14676\,
            in3 => \N__14772\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIRHJAF_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__19434\,
            in1 => \N__23349\,
            in2 => \N__14667\,
            in3 => \N__16251\,
            lcout => \Lab_UT.scctrl.next_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_0_RNIJFLD2_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__22191\,
            in1 => \N__22460\,
            in2 => \N__19730\,
            in3 => \N__22029\,
            lcout => \Lab_UT.scctrl.N_415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNIBUL06_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21501\,
            in1 => \N__21377\,
            in2 => \N__20662\,
            in3 => \N__22190\,
            lcout => \Lab_UT.scctrl.N_401_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_4_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20651\,
            in1 => \N__22641\,
            in2 => \N__21409\,
            in3 => \N__21502\,
            lcout => \Lab_UT.scctrl.G_24_i_a7_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_8_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100011"
        )
    port map (
            in0 => \N__22028\,
            in1 => \N__18282\,
            in2 => \N__19945\,
            in3 => \N__23108\,
            lcout => \Lab_UT.scctrl.next_state_rst_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIN79O4_0_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23348\,
            in1 => \N__21390\,
            in2 => \N__18954\,
            in3 => \N__21500\,
            lcout => \Lab_UT.scctrl.G_15_0_a10_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_9_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100001111"
        )
    port map (
            in0 => \N__21499\,
            in1 => \N__16212\,
            in2 => \N__19156\,
            in3 => \N__23117\,
            lcout => \Lab_UT.scctrl.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNIKFLC4_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111111111"
        )
    port map (
            in0 => \N__21388\,
            in1 => \N__22037\,
            in2 => \N__19941\,
            in3 => \N__21498\,
            lcout => \Lab_UT.scctrl.g0_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_2_rep1_RNI4P8F2_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__20451\,
            in1 => \N__16211\,
            in2 => \_gnd_net_\,
            in3 => \N__22175\,
            lcout => \Lab_UT.scctrl.g0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_3_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22177\,
            in1 => \N__14762\,
            in2 => \N__19157\,
            in3 => \N__16210\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_419_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__19492\,
            in1 => \N__23463\,
            in2 => \N__14745\,
            in3 => \N__15225\,
            lcout => \Lab_UT.scctrl.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_6_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__21389\,
            in1 => \N__20647\,
            in2 => \N__14730\,
            in3 => \N__15450\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_2_RNO_2_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__15234\,
            in1 => \N__19144\,
            in2 => \N__15228\,
            in3 => \N__23118\,
            lcout => \Lab_UT.scctrl.g0_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__22176\,
            in1 => \N__22792\,
            in2 => \N__22461\,
            in3 => \N__22036\,
            lcout => \Lab_UT.scctrl.N_418_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_3_RNI7ARC1_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14852\,
            in1 => \N__16560\,
            in2 => \N__14949\,
            in3 => \N__17890\,
            lcout => \Lab_UT.scctrl.N_444_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_3_RNI7ARC1_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14941\,
            in1 => \N__16559\,
            in2 => \N__17898\,
            in3 => \N__14851\,
            lcout => \Lab_UT.scctrl.N_444_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_7_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16208\,
            in1 => \N__15195\,
            in2 => \N__20456\,
            in3 => \N__15129\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_24_i_a6_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011000"
        )
    port map (
            in0 => \N__22236\,
            in1 => \N__22826\,
            in2 => \N__14964\,
            in3 => \N__15243\,
            lcout => \Lab_UT.scctrl.G_24_i_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_4_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16209\,
            in1 => \N__17891\,
            in2 => \N__18087\,
            in3 => \N__22235\,
            lcout => \Lab_UT.scctrl.G_24_i_a6_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_5_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__16561\,
            in1 => \N__14961\,
            in2 => \N__14948\,
            in3 => \N__14853\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__14820\,
            in1 => \N__14814\,
            in2 => \N__14808\,
            in3 => \N__15318\,
            lcout => \Lab_UT.scctrl.next_state_rst_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_2_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111101"
        )
    port map (
            in0 => \N__23607\,
            in1 => \N__16029\,
            in2 => \N__18085\,
            in3 => \N__23119\,
            lcout => \Lab_UT.scctrl.G_24_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__15311\,
            in1 => \N__15291\,
            in2 => \N__18439\,
            in3 => \N__15264\,
            lcout => \Lab_UT.scctrl.next_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21081\,
            ce => \N__20899\,
            sr => \N__20857\
        );

    \Lab_UT.scctrl.state_ret_RNIKML91_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__16013\,
            in1 => \N__18420\,
            in2 => \_gnd_net_\,
            in3 => \N__22057\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_170_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_RNIK5UKH_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15498\,
            in1 => \_gnd_net_\,
            in2 => \N__15246\,
            in3 => \N__17457\,
            lcout => \Lab_UT.state_ret_RNIK5UKH_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_12_RNIUVHQG_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__17952\,
            in1 => \N__19814\,
            in2 => \N__16017\,
            in3 => \N__15499\,
            lcout => \Lab_UT.state_ret_12_RNIUVHQG_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_8_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22442\,
            in2 => \_gnd_net_\,
            in3 => \N__22053\,
            lcout => \Lab_UT.scctrl.G_24_i_o6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_12_RNI2D6E_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19813\,
            in1 => \N__19158\,
            in2 => \_gnd_net_\,
            in3 => \N__22802\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_17_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_12_RNI2SEPG_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15497\,
            in1 => \_gnd_net_\,
            in2 => \N__15237\,
            in3 => \N__17358\,
            lcout => \Lab_UT.state_ret_12_RNI2SEPG_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI2IGHH_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18488\,
            in1 => \N__15990\,
            in2 => \_gnd_net_\,
            in3 => \N__15496\,
            lcout => \Lab_UT.state_1_RNI2IGHH_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIOII81_2_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19154\,
            in1 => \N__22823\,
            in2 => \N__18440\,
            in3 => \N__22055\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_20_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIO1RJH_2_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__17549\,
            in1 => \_gnd_net_\,
            in2 => \N__15537\,
            in3 => \N__15494\,
            lcout => \Lab_UT.state_1_RNIO1RJH_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNILCGA1_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111110001"
        )
    port map (
            in0 => \N__19153\,
            in1 => \N__22822\,
            in2 => \N__20691\,
            in3 => \N__16012\,
            lcout => \Lab_UT.scctrl.N_277\,
            ltout => \Lab_UT.scctrl.N_277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNIR2443_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__22976\,
            in1 => \N__15510\,
            in2 => \N__15528\,
            in3 => \N__18906\,
            lcout => \N_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_RNIVRBS_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18427\,
            in1 => \N__22825\,
            in2 => \_gnd_net_\,
            in3 => \N__22056\,
            lcout => \Lab_UT.scctrl.N_355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNI2KLS_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__22824\,
            in1 => \N__20690\,
            in2 => \_gnd_net_\,
            in3 => \N__19155\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_27_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNI23U7H_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15495\,
            in1 => \_gnd_net_\,
            in2 => \N__15465\,
            in3 => \N__17508\,
            lcout => \Lab_UT.state_1_ret_3_RNI23U7H_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_3_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110011"
        )
    port map (
            in0 => \N__23488\,
            in1 => \N__15462\,
            in2 => \N__15327\,
            in3 => \N__19340\,
            lcout => \Lab_UT.scctrl.G_18_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_2_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__15567\,
            in1 => \N__15588\,
            in2 => \N__23708\,
            in3 => \N__23494\,
            lcout => \Lab_UT.scctrl.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20826\
        );

    \Lab_UT.scctrl.state_1_fast_2_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__23491\,
            in1 => \N__23705\,
            in2 => \N__15597\,
            in3 => \N__15570\,
            lcout => \Lab_UT.scctrl.state_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20826\
        );

    \Lab_UT.scctrl.state_1_2_rep1_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__15568\,
            in1 => \N__15589\,
            in2 => \N__23709\,
            in3 => \N__23495\,
            lcout => \Lab_UT.scctrl.state_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20826\
        );

    \Lab_UT.scctrl.state_ret_0_RNI1ME69_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__22296\,
            in1 => \N__15654\,
            in2 => \N__15711\,
            in3 => \N__21522\,
            lcout => \Lab_UT.scctrl.g1_2_0\,
            ltout => \Lab_UT.scctrl.g1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNI3K1MC_2_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23697\,
            in1 => \N__15587\,
            in2 => \N__15648\,
            in3 => \N__23489\,
            lcout => \Lab_UT.scctrl.next_stateZ0Z_2\,
            ltout => \Lab_UT.scctrl.next_stateZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001111110111111"
        )
    port map (
            in0 => \N__23492\,
            in1 => \N__19530\,
            in2 => \N__15645\,
            in3 => \N__15641\,
            lcout => \Lab_UT.scctrl.N_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20826\
        );

    \Lab_UT.scctrl.state_ret_1_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__15642\,
            in1 => \N__23493\,
            in2 => \N__19536\,
            in3 => \N__15613\,
            lcout => \Lab_UT.scctrl.N_296_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20826\
        );

    \Lab_UT.scctrl.state_1_2_rep2_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__23490\,
            in1 => \N__23704\,
            in2 => \N__15596\,
            in3 => \N__15569\,
            lcout => \Lab_UT.scctrl.state_2_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21143\,
            ce => 'H',
            sr => \N__20826\
        );

    \Lab_UT.scctrl.state_1_ret_5_RNO_4_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100011"
        )
    port map (
            in0 => \N__21996\,
            in1 => \N__18230\,
            in2 => \N__19944\,
            in3 => \N__23186\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_5_RNO_2_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__18432\,
            in1 => \N__15698\,
            in2 => \N__15555\,
            in3 => \N__15552\,
            lcout => \Lab_UT.scctrl.g0_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNO_5_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100011"
        )
    port map (
            in0 => \N__21993\,
            in1 => \N__18225\,
            in2 => \N__19942\,
            in3 => \N__23183\,
            lcout => \Lab_UT.scctrl.next_state_rst_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNO_5_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101011"
        )
    port map (
            in0 => \N__23185\,
            in1 => \N__19926\,
            in2 => \N__18259\,
            in3 => \N__21997\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_4_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNO_2_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__15697\,
            in1 => \N__18431\,
            in2 => \N__15720\,
            in3 => \N__15717\,
            lcout => \Lab_UT.scctrl.g0_2_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_2_rep2_RNI2S7K1_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__21315\,
            in1 => \N__21994\,
            in2 => \N__18054\,
            in3 => \N__22918\,
            lcout => \Lab_UT.scctrl.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNI1HVT2_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100011"
        )
    port map (
            in0 => \N__21995\,
            in1 => \N__18226\,
            in2 => \N__19943\,
            in3 => \N__23184\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_RNI227Q7_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__18430\,
            in1 => \N__15696\,
            in2 => \N__15672\,
            in3 => \N__15669\,
            lcout => \Lab_UT.scctrl.g0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIB2MFC_3_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__19242\,
            in1 => \N__19521\,
            in2 => \N__23498\,
            in3 => \N__15787\,
            lcout => \Lab_UT.scctrl.next_state_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_fast_3_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__15790\,
            in1 => \N__23426\,
            in2 => \N__19535\,
            in3 => \N__19245\,
            lcout => \Lab_UT.scctrl.state_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => 'H',
            sr => \N__20823\
        );

    \Lab_UT.scctrl.state_2_3_rep1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__19244\,
            in1 => \N__19525\,
            in2 => \N__23499\,
            in3 => \N__15789\,
            lcout => \Lab_UT.scctrl.state_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => 'H',
            sr => \N__20823\
        );

    \Lab_UT.scctrl.state_2_3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__15788\,
            in1 => \N__23425\,
            in2 => \N__19534\,
            in3 => \N__19243\,
            lcout => \Lab_UT.scctrl.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => 'H',
            sr => \N__20823\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNO_2_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__22290\,
            in1 => \N__22400\,
            in2 => \N__22044\,
            in3 => \N__22737\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_418_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNO_0_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__19520\,
            in1 => \N__23421\,
            in2 => \N__15807\,
            in3 => \N__19241\,
            lcout => \Lab_UT.scctrl.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_6_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111001101010011"
        )
    port map (
            in0 => \N__19246\,
            in1 => \N__19529\,
            in2 => \N__23500\,
            in3 => \N__15791\,
            lcout => \Lab_UT.scctrl.state_i_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21130\,
            ce => 'H',
            sr => \N__20823\
        );

    \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100010"
        )
    port map (
            in0 => \N__22736\,
            in1 => \N__21989\,
            in2 => \N__22440\,
            in3 => \N__22289\,
            lcout => \Lab_UT.scctrl.N_418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011000110111011"
        )
    port map (
            in0 => \N__23433\,
            in1 => \N__23691\,
            in2 => \N__15765\,
            in3 => \N__18113\,
            lcout => \Lab_UT.scctrl.state_i_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21125\,
            ce => 'H',
            sr => \N__20822\
        );

    \Lab_UT.scctrl.state_ret_0_fast_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110100001111"
        )
    port map (
            in0 => \N__18114\,
            in1 => \N__15764\,
            in2 => \N__23707\,
            in3 => \N__23434\,
            lcout => \Lab_UT.scctrl.state_ret_0_fastZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21125\,
            ce => 'H',
            sr => \N__20822\
        );

    \Lab_UT.scctrl.state_ret_0_RNIKR11_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23394\,
            in2 => \_gnd_net_\,
            in3 => \N__19669\,
            lcout => \Lab_UT.scctrl.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_11_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__15742\,
            in1 => \_gnd_net_\,
            in2 => \N__23487\,
            in3 => \N__22769\,
            lcout => \Lab_UT.scctrl.G_18_i_a9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_10_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16279\,
            in2 => \_gnd_net_\,
            in3 => \N__15741\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.state_ret_4_RNOZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNO_6_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111110101"
        )
    port map (
            in0 => \N__20520\,
            in1 => \N__20641\,
            in2 => \N__16032\,
            in3 => \N__21364\,
            lcout => \Lab_UT.scctrl.state_ret_4_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_0_RNIJOQD_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19670\,
            in2 => \_gnd_net_\,
            in3 => \N__22888\,
            lcout => \Lab_UT.scctrl.N_295\,
            ltout => \Lab_UT.scctrl.N_295_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI23861_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21365\,
            in2 => \N__15993\,
            in3 => \N__21960\,
            lcout => \Lab_UT.scctrl.N_40_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15978\,
            in1 => \N__15924\,
            in2 => \_gnd_net_\,
            in3 => \N__15900\,
            lcout => \Lab_UT.scctrl.next_state_rst_0_3_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_2_rep1_RNIJJLN1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__21974\,
            in1 => \N__20452\,
            in2 => \N__16575\,
            in3 => \N__16104\,
            lcout => \Lab_UT.scctrl.N_408\,
            ltout => \Lab_UT.scctrl.N_408_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_16_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__16040\,
            in1 => \N__16218\,
            in2 => \N__15837\,
            in3 => \N__23179\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_i_a8_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_9_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__21975\,
            in1 => \N__16328\,
            in2 => \N__15834\,
            in3 => \N__19976\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_12_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_2_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__19247\,
            in1 => \N__15831\,
            in2 => \N__15819\,
            in3 => \N__19268\,
            lcout => \Lab_UT.scctrl.N_13_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNO_0_1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__23180\,
            in1 => \N__18147\,
            in2 => \N__15816\,
            in3 => \N__16041\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__16329\,
            in1 => \N__19977\,
            in2 => \N__16320\,
            in3 => \N__21976\,
            lcout => \Lab_UT.scctrl.next_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21119\,
            ce => \N__20901\,
            sr => \N__20846\
        );

    \Lab_UT.scctrl.state_2_fast_RNI7HMP_3_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__16317\,
            in1 => \N__18898\,
            in2 => \_gnd_net_\,
            in3 => \N__16281\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_5_RNI7FV82_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__16163\,
            in1 => \N__16192\,
            in2 => \N__16257\,
            in3 => \N__16230\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_1_RNIGQ5R4_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__18247\,
            in1 => \N__16224\,
            in2 => \N__16254\,
            in3 => \N__23162\,
            lcout => \Lab_UT.scctrl.g0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_fast_RNIFRSV_2_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__20375\,
            in1 => \N__21965\,
            in2 => \N__16164\,
            in3 => \N__16245\,
            lcout => \Lab_UT.scctrl.N_408_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_rep1_RNI9FBG_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19907\,
            in2 => \_gnd_net_\,
            in3 => \N__20512\,
            lcout => \Lab_UT.scctrl.g2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_19_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011111"
        )
    port map (
            in0 => \N__20513\,
            in1 => \_gnd_net_\,
            in2 => \N__19934\,
            in3 => \N__18246\,
            lcout => \Lab_UT.scctrl.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_5_RNIH2CF_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16191\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16162\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNIJOFP1_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__18899\,
            in1 => \N__23573\,
            in2 => \N__16044\,
            in3 => \N__19596\,
            lcout => \Lab_UT.scctrl.next_state_rst_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__19749\,
            in1 => \N__16380\,
            in2 => \N__22593\,
            in3 => \N__16467\,
            lcout => \Lab_UT.scctrl.nibbleInZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21105\,
            ce => \N__16497\,
            sr => \N__16371\
        );

    \Lab_UT.scctrl.shifter_ret_7_RNIQ5993_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__21972\,
            in1 => \N__22449\,
            in2 => \N__16485\,
            in3 => \N__22196\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_69_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNI6DT75_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000100010"
        )
    port map (
            in0 => \N__21570\,
            in1 => \N__16466\,
            in2 => \N__16458\,
            in3 => \N__19748\,
            lcout => \Lab_UT.sccDnibble1En\,
            ltout => \Lab_UT.sccDnibble1En_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_esr_RNO_2_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16455\,
            in3 => \N__16452\,
            lcout => \Lab_UT.scdp.u0.sccDnibble1En_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_7_RNIEAT93_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__22198\,
            in1 => \N__16395\,
            in2 => \N__22463\,
            in3 => \N__21973\,
            lcout => \Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93\,
            ltout => \Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16374\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scctrl.N_69_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_10_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__21971\,
            in1 => \N__22450\,
            in2 => \N__19031\,
            in3 => \N__22197\,
            lcout => \Lab_UT.scctrl.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIDAFVC_3_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__19620\,
            in1 => \N__23196\,
            in2 => \N__22977\,
            in3 => \N__16671\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_9_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIN96CP1_3_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000010000"
        )
    port map (
            in0 => \N__16358\,
            in1 => \N__16716\,
            in2 => \N__16332\,
            in3 => \N__20017\,
            lcout => \Lab_UT.scctrl.next_state_RNIN96CP1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.shifter_ret_3_RNIV6006_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__16755\,
            in1 => \N__16743\,
            in2 => \_gnd_net_\,
            in3 => \N__16730\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g1_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNICEBUC_3_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__23454\,
            in1 => \N__19518\,
            in2 => \N__16719\,
            in3 => \N__16677\,
            lcout => \Lab_UT.scctrl.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI91NK6_2_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__19103\,
            in1 => \N__16710\,
            in2 => \N__16704\,
            in3 => \N__23195\,
            lcout => \Lab_UT.scctrl.g0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIDJ6B1_2_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__20313\,
            in1 => \N__19104\,
            in2 => \N__18429\,
            in3 => \N__22815\,
            lcout => \Lab_UT.scctrl.g0_9_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_3_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__21537\,
            in1 => \N__16661\,
            in2 => \N__17913\,
            in3 => \N__17893\,
            lcout => \Lab_UT.scdp.byteToDecrypt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21093\,
            ce => 'H',
            sr => \N__20825\
        );

    \Lab_UT.scdp.a2b.val_i_0_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__17055\,
            in1 => \N__16643\,
            in2 => \N__17206\,
            in3 => \N__17074\,
            lcout => \Lab_UT.scdp.val_i_0_0\,
            ltout => \Lab_UT.scdp.val_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.rxdataD.q_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16647\,
            in3 => \N__17276\,
            lcout => \Lab_UT.scdp.binValD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21093\,
            ce => 'H',
            sr => \N__20825\
        );

    \Lab_UT.scdp.a2b.val_i_a2_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__16644\,
            in1 => \N__17195\,
            in2 => \N__16581\,
            in3 => \N__17075\,
            lcout => \Lab_UT.scdp.N_378\,
            ltout => \Lab_UT.scdp.N_378_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__17291\,
            in1 => \N__17306\,
            in2 => \N__17313\,
            in3 => \N__16951\,
            lcout => \Lab_UT.scdp.byteToDecrypt_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21093\,
            ce => 'H',
            sr => \N__20825\
        );

    \Lab_UT.scdp.u1.q_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__17292\,
            in1 => \N__17251\,
            in2 => \N__17280\,
            in3 => \N__21536\,
            lcout => \Lab_UT.scdp.u1.byteToDecryptZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21093\,
            ce => 'H',
            sr => \N__20825\
        );

    \Lab_UT.scdp.a2b.shifter_ret_RNIJ2EC2_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__17232\,
            in1 => \N__17191\,
            in2 => \N__17076\,
            in3 => \N__17054\,
            lcout => \Lab_UT.scdp.val_0_tz_3\,
            ltout => \Lab_UT.scdp.val_0_tz_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_3_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__16952\,
            in1 => \N__16926\,
            in2 => \N__16932\,
            in3 => \N__17892\,
            lcout => \Lab_UT.scdp.byteToDecrypt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21093\,
            ce => 'H',
            sr => \N__20825\
        );

    \Lab_UT.scdp.k2l.q_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17600\,
            in1 => \N__18685\,
            in2 => \N__16907\,
            in3 => \N__17453\,
            lcout => \Lab_UT.scdp.key2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21088\,
            ce => 'H',
            sr => \N__20828\
        );

    \Lab_UT.scdp.k2l.q_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__17454\,
            in1 => \N__18676\,
            in2 => \N__16886\,
            in3 => \N__17408\,
            lcout => \Lab_UT.scdp.key2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21088\,
            ce => 'H',
            sr => \N__20828\
        );

    \Lab_UT.scdp.k3l.q_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17601\,
            in1 => \N__18686\,
            in2 => \N__16868\,
            in3 => \N__17948\,
            lcout => \Lab_UT.scdp.key3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21088\,
            ce => 'H',
            sr => \N__20828\
        );

    \Lab_UT.scdp.k3l.q_1_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__17949\,
            in1 => \N__18677\,
            in2 => \N__16844\,
            in3 => \N__17409\,
            lcout => \Lab_UT.scdp.key3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21088\,
            ce => 'H',
            sr => \N__20828\
        );

    \Lab_UT.scdp.k3l.q_2_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18675\,
            in1 => \N__16826\,
            in2 => \N__16772\,
            in3 => \N__17950\,
            lcout => \Lab_UT.scdp.key3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21088\,
            ce => 'H',
            sr => \N__20828\
        );

    \Lab_UT.scdp.k3l.q_3_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__17951\,
            in1 => \N__18678\,
            in2 => \N__17930\,
            in3 => \N__18517\,
            lcout => \Lab_UT.scdp.key3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21088\,
            ce => 'H',
            sr => \N__20828\
        );

    \Lab_UT.scdp.rxdataD.q_3_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17909\,
            in2 => \_gnd_net_\,
            in3 => \N__17886\,
            lcout => \Lab_UT.scdp.binValD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21088\,
            ce => 'H',
            sr => \N__20828\
        );

    \buart.Z_rx.hh_RNIJ3K62_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__17792\,
            in1 => \N__17763\,
            in2 => \_gnd_net_\,
            in3 => \N__17734\,
            lcout => \buart.Z_rx.startbit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.k0l.q_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18679\,
            in1 => \N__17615\,
            in2 => \N__17573\,
            in3 => \N__17544\,
            lcout => \Lab_UT.scdp.key0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21082\,
            ce => 'H',
            sr => \N__20829\
        );

    \Lab_UT.scdp.k0l.q_1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__17545\,
            in1 => \N__17393\,
            in2 => \N__17525\,
            in3 => \N__18682\,
            lcout => \Lab_UT.scdp.key0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21082\,
            ce => 'H',
            sr => \N__20829\
        );

    \Lab_UT.scdp.k1h.q_1_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18683\,
            in1 => \N__17394\,
            in2 => \N__17474\,
            in3 => \N__17504\,
            lcout => \Lab_UT.scdp.key1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21082\,
            ce => 'H',
            sr => \N__20829\
        );

    \Lab_UT.scdp.k2l.q_3_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18681\,
            in1 => \N__18516\,
            in2 => \N__17426\,
            in3 => \N__17456\,
            lcout => \Lab_UT.scdp.key2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21082\,
            ce => 'H',
            sr => \N__20829\
        );

    \Lab_UT.scdp.k1l.q_1_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18684\,
            in1 => \N__17395\,
            in2 => \N__17330\,
            in3 => \N__17357\,
            lcout => \Lab_UT.scdp.key1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21082\,
            ce => 'H',
            sr => \N__20829\
        );

    \Lab_UT.scdp.k2h.q_3_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__18680\,
            in1 => \N__18515\,
            in2 => \N__18458\,
            in3 => \N__18484\,
            lcout => \Lab_UT.scdp.key2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21082\,
            ce => 'H',
            sr => \N__20829\
        );

    \Lab_UT.scctrl.next_state_RNO_1_1_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__18428\,
            in1 => \N__19930\,
            in2 => \_gnd_net_\,
            in3 => \N__18276\,
            lcout => \Lab_UT.scctrl.next_state_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_2_rep2_RNIB7181_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22963\,
            in1 => \N__21961\,
            in2 => \_gnd_net_\,
            in3 => \N__18066\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIE6PO6_0_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21416\,
            in1 => \N__22288\,
            in2 => \N__18132\,
            in3 => \N__21521\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIMNKBA_3_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000100"
        )
    port map (
            in0 => \N__22965\,
            in1 => \N__18129\,
            in2 => \N__18117\,
            in3 => \N__23188\,
            lcout => \Lab_UT.scctrl.next_state_rst_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_0_RNO_5_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__18067\,
            in1 => \_gnd_net_\,
            in2 => \N__22035\,
            in3 => \N__22964\,
            lcout => \Lab_UT.scctrl.N_319_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_10_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19599\,
            in1 => \N__18072\,
            in2 => \_gnd_net_\,
            in3 => \N__21818\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_5_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21403\,
            in1 => \N__23509\,
            in2 => \N__17955\,
            in3 => \N__21520\,
            lcout => \Lab_UT.scctrl.G_18_i_a9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_4_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__19164\,
            in1 => \N__23182\,
            in2 => \N__23523\,
            in3 => \N__22957\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_18_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_0_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__18978\,
            in1 => \N__18972\,
            in2 => \N__18960\,
            in3 => \N__22291\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_18_i_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19188\,
            in1 => \N__19215\,
            in2 => \N__18957\,
            in3 => \N__20055\,
            lcout => \Lab_UT.scctrl.N_398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_10_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21817\,
            in1 => \N__20434\,
            in2 => \_gnd_net_\,
            in3 => \N__19598\,
            lcout => \Lab_UT.scctrl.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNICEV81_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__19935\,
            in1 => \N__21402\,
            in2 => \N__21949\,
            in3 => \N__20179\,
            lcout => \Lab_UT.scctrl.state_1_ret_1_RNICEVZ0Z81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_2_rep1_RNI8F771_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21816\,
            in1 => \N__20433\,
            in2 => \_gnd_net_\,
            in3 => \N__19597\,
            lcout => \Lab_UT.scctrl.N_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_RNO_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__23506\,
            in1 => \N__18936\,
            in2 => \N__20288\,
            in3 => \N__18924\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_4_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20181\,
            in2 => \N__18909\,
            in3 => \N__20053\,
            lcout => \Lab_UT.scctrl.N_260_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21131\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_1_0_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__18861\,
            in1 => \N__22830\,
            in2 => \N__18831\,
            in3 => \N__18812\,
            lcout => \Lab_UT.scctrl.g0_1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20180\,
            in2 => \_gnd_net_\,
            in3 => \N__20052\,
            lcout => \Lab_UT.scctrl.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21131\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_2_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011110101111"
        )
    port map (
            in0 => \N__23505\,
            in1 => \N__19272\,
            in2 => \N__20289\,
            in3 => \N__19251\,
            lcout => \Lab_UT.scctrl.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_6_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23672\,
            in2 => \_gnd_net_\,
            in3 => \N__19519\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__19209\,
            in1 => \N__23504\,
            in2 => \N__19191\,
            in3 => \N__19390\,
            lcout => \Lab_UT.scctrl.N_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNO_9_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__22436\,
            in1 => \N__21872\,
            in2 => \N__19179\,
            in3 => \N__22287\,
            lcout => \Lab_UT.scctrl.N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_11_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__22258\,
            in1 => \N__19133\,
            in2 => \N__19035\,
            in3 => \N__23178\,
            lcout => \Lab_UT.scctrl.N_21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_14_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__22432\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21854\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_10_i_o7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_7_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__22259\,
            in1 => \N__19727\,
            in2 => \N__18993\,
            in3 => \N__23508\,
            lcout => \Lab_UT.scctrl.N_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_0_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__21204\,
            in1 => \N__18990\,
            in2 => \N__22592\,
            in3 => \N__22260\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_24_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__22637\,
            in1 => \N__22470\,
            in2 => \N__19761\,
            in3 => \N__19758\,
            lcout => \Lab_UT.scctrl.rst_retZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_0_RNIJFLD2_2_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__21858\,
            in1 => \N__19726\,
            in2 => \N__22458\,
            in3 => \N__22256\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_0_RNIUTK59_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__22257\,
            in1 => \N__19542\,
            in2 => \N__19632\,
            in3 => \N__19629\,
            lcout => \Lab_UT.scctrl.g0_9_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_2_rep1_RNIV3EJ1_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__21404\,
            in1 => \N__19607\,
            in2 => \N__20457\,
            in3 => \N__21853\,
            lcout => \Lab_UT.scctrl.g0_9_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNIU5BF_4_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22582\,
            in2 => \_gnd_net_\,
            in3 => \N__23443\,
            lcout => \N_21_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_18_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__19494\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20250\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.m90_i_o6_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_13_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__19433\,
            in1 => \N__22583\,
            in2 => \N__19410\,
            in3 => \N__23444\,
            lcout => \Lab_UT.scctrl.N_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_5_RNO_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19407\,
            in1 => \N__19391\,
            in2 => \_gnd_net_\,
            in3 => \N__19341\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_5_RNO_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__20252\,
            in1 => \N__23448\,
            in2 => \N__19287\,
            in3 => \N__19284\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_5_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001010"
        )
    port map (
            in0 => \N__22584\,
            in1 => \N__20140\,
            in2 => \N__20331\,
            in3 => \N__20054\,
            lcout => \Lab_UT.scctrl.N_356_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_4_RNIDMQE_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__23604\,
            in1 => \N__20139\,
            in2 => \_gnd_net_\,
            in3 => \N__23442\,
            lcout => \Lab_UT.scctrl.g0_9_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNO_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__20301\,
            in1 => \N__20251\,
            in2 => \N__23502\,
            in3 => \N__20196\,
            lcout => \Lab_UT.scctrl.next_state_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_3_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__20182\,
            in1 => \N__20061\,
            in2 => \_gnd_net_\,
            in3 => \N__20045\,
            lcout => \Lab_UT.scctrl.N_260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIFADO_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21413\,
            in2 => \_gnd_net_\,
            in3 => \N__21928\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_1_i_i_a2_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_ret_1_RNI4KSC6_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111111"
        )
    port map (
            in0 => \N__19946\,
            in1 => \N__22194\,
            in2 => \N__19980\,
            in3 => \N__21518\,
            lcout => \Lab_UT.scctrl.next_state_rst_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNIP7S81_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__19956\,
            in1 => \N__21414\,
            in2 => \N__22030\,
            in3 => \N__19947\,
            lcout => \N_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_RNIOCR32_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22428\,
            in1 => \N__19815\,
            in2 => \N__19788\,
            in3 => \N__22193\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_72_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_RNI4RQC3_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__21187\,
            in1 => \N__19770\,
            in2 => \N__21627\,
            in3 => \N__21608\,
            lcout => \Lab_UT.state_ret_11_RNI4RQC3_0\,
            ltout => \Lab_UT.state_ret_11_RNI4RQC3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNIP7S81_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21597\,
            in3 => \N__21561\,
            lcout => \Lab_UT.sccDnibble2En\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_3_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21519\,
            in1 => \N__21415\,
            in2 => \N__21219\,
            in3 => \N__23513\,
            lcout => \Lab_UT.scctrl.G_10_i_a7_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_2_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21188\,
            lcout => \Lab_UT.scctrl.next_state_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21107\,
            ce => \N__20892\,
            sr => \N__20858\
        );

    \Lab_UT.scctrl.state_1_ret_3_RNIJURV_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__20686\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20663\,
            lcout => \N_55_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_17_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__20524\,
            in1 => \N__23503\,
            in2 => \N__20447\,
            in3 => \N__22821\,
            lcout => \Lab_UT.scctrl.N_13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_11_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110111"
        )
    port map (
            in0 => \N__23440\,
            in1 => \N__23606\,
            in2 => \N__23695\,
            in3 => \N__20391\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_10_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_5_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__22962\,
            in1 => \N__23198\,
            in2 => \N__20385\,
            in3 => \N__23441\,
            lcout => \Lab_UT.scctrl.G_10_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_fast_RNIM0M4_2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__20382\,
            in1 => \N__22788\,
            in2 => \N__23501\,
            in3 => \N__20358\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIMPVR_2_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110111"
        )
    port map (
            in0 => \N__23668\,
            in1 => \N__23605\,
            in2 => \N__23532\,
            in3 => \N__23438\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_15_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIKG4B3_3_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__23439\,
            in1 => \N__23181\,
            in2 => \N__22980\,
            in3 => \N__22961\,
            lcout => \Lab_UT.scctrl.G_15_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_6_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__22789\,
            in1 => \N__22636\,
            in2 => \N__22617\,
            in3 => \N__21735\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_24_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_1_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__22608\,
            in1 => \N__22602\,
            in2 => \N__22596\,
            in3 => \N__22585\,
            lcout => \Lab_UT.scctrl.G_24_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.rst_ret_RNO_12_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__22459\,
            in1 => \N__22195\,
            in2 => \_gnd_net_\,
            in3 => \N__21948\,
            lcout => \Lab_UT.scctrl.N_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNICOE1_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21722\,
            lcout => \N_245_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
