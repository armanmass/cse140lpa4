-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Jun 3 2019 04:04:59

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__23195\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \latticehx1k_pll_inst.clk\ : std_logic;
signal clk_in_c : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.N_41_i\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal \uart_RXD\ : std_logic;
signal \bfn_2_5_0_\ : std_logic;
signal \buart.Z_tx.counter_RNIVE1P1_1\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_0\ : std_logic;
signal \buart.Z_tx.counter_RNIVE1P1_0_1\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_1\ : std_logic;
signal \buart.Z_tx.un1_bitcount_axb_3\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_2\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \ufifo.fifo.fifo_txdata_2\ : std_logic;
signal \ufifo.fifo.fifo_txdata_1\ : std_logic;
signal \ufifo.sb_ram512x8_inst_RNIKRN11_cascade_\ : std_logic;
signal \ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0\ : std_logic;
signal utb_txdata_1 : std_logic;
signal \ufifo.fifo.fifo_txdata_0\ : std_logic;
signal \ufifo.fifo.fifo_txdata_6\ : std_logic;
signal \ufifo.fifo.fifo_txdata_5\ : std_logic;
signal ufifo_utb_txdata_m0_5 : std_logic;
signal \ufifo.fifo.fifo_txdata_7\ : std_logic;
signal ufifo_utb_txdata_m0_7 : std_logic;
signal ufifo_utb_txdata_m0_6 : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal \ufifo.un4_rxDataValidNoEscZ0Z_1_cascade_\ : std_logic;
signal \ufifo.rxDataValidNoEscZ0\ : std_logic;
signal \ufifo.fifo.fifo_txdata_3\ : std_logic;
signal \ufifo.fifo.fifo_txdata_4\ : std_logic;
signal \ufifo.utb_txdata_m0_0\ : std_logic;
signal utb_txdata_0 : std_logic;
signal \Lab_UT_dk_de_cr_2_reti\ : std_logic;
signal ufifo_utb_txdata_m0_3 : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal ufifo_utb_txdata_m0_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_7\ : std_logic;
signal \Lab_UT.scdp.u2.byteToEncrypt_0\ : std_logic;
signal \bfn_4_1_0_\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_0\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_1\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_2\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_3\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_4\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_5\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_6\ : std_logic;
signal \ufifo.fifo.un1_rdaddr_cry_7\ : std_logic;
signal \bfn_4_2_0_\ : std_logic;
signal \bfn_4_3_0_\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_0\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_1\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_2\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_3\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_4\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_5\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_6\ : std_logic;
signal \ufifo.fifo.un1_wraddr_cry_7\ : std_logic;
signal \bfn_4_4_0_\ : std_logic;
signal \resetGen.un12_ci_cascade_\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_6\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_7\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_7\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_6\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_0\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_8\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_8\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_0\ : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \Lab_UT.scdp.q_RNI56C1D_0_cascade_\ : std_logic;
signal \ufifo.txdataDZ0Z_0\ : std_logic;
signal \ufifo.txdataDZ0Z_6\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \resetGen.reset_count_2_0_4_cascade_\ : std_logic;
signal \resetGen.un12_ci\ : std_logic;
signal \resetGen.un23_ci\ : std_logic;
signal \resetGen.escKeyZ0\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \Lab_UT.scdp.msBitsi.q_esr_RNIF1M8Z0Z_6\ : std_logic;
signal \Lab_UT.scdp.msBitsi.q_esr_RNIQQ8EZ0Z_0\ : std_logic;
signal \resetGen.escKey_0Z0Z_0\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsD_6\ : std_logic;
signal \Lab_UT.scdp.u2.byteToEncryptZ0Z_5\ : std_logic;
signal \Lab_UT.scdp.d2eData_5_cascade_\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_6\ : std_logic;
signal \Lab_UT.scdp.N_52_cascade_\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsDZ0Z_0\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_4\ : std_logic;
signal \Lab_UT.scdp.b2a0.N_55\ : std_logic;
signal \Lab_UT.scdp.d2eData_5\ : std_logic;
signal \Lab_UT.scdp.b2a0.N_55_cascade_\ : std_logic;
signal \Lab_UT.scdp.a2b.val_0_0Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_6\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_6_cascade_\ : std_logic;
signal \Lab_UT.scdp.u0.byteToDecrypt_6\ : std_logic;
signal \ufifo.sb_ram512x8_inst_RNILSN11\ : std_logic;
signal \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0_cascade_\ : std_logic;
signal ufifo_utb_txdata_sm0_0 : std_logic;
signal utb_txdata_2 : std_logic;
signal \ufifo.txdataDZ0Z_1\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsD_1\ : std_logic;
signal \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8Z0Z_1\ : std_logic;
signal \ufifo.txdataDZ0Z_5\ : std_logic;
signal \Lab_UT.scdp.u2.sccEldByte_0\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsD_2\ : std_logic;
signal \Lab_UT.scdp.msBitsi.L4_tx_data_ns_1_2_cascade_\ : std_logic;
signal \ufifo.txdataDZ0Z_2\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_1_cascade_\ : std_logic;
signal \Lab_UT.scdp.q_RNIABC1D_1\ : std_logic;
signal \Lab_UT.scdp.u2.byteToEncrypt_1\ : std_logic;
signal \Lab_UT.scdp.d2eData_1_cascade_\ : std_logic;
signal \Lab_UT.scdp.lsBits_6_cascade_\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_1\ : std_logic;
signal \Lab_UT.scdp.lsBitsi.lsBitsD_3\ : std_logic;
signal \Lab_UT.scdp.byteToEncrypt_3\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_6\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_2_cascade_\ : std_logic;
signal \Lab_UT.scdp.u2.byteToEncrypt_2\ : std_logic;
signal \Lab_UT.scdp.d2eData_2\ : std_logic;
signal \Lab_UT.scdp.d2eData_1\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_2\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_1\ : std_logic;
signal \Lab_UT.scdp.pinst0.un12_pValidZ0Z_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.un12_pValid_cascade_\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_0\ : std_logic;
signal \Lab_UT.scdp.un12_pValid\ : std_logic;
signal \Lab_UT.scdp.e2dData_6\ : std_logic;
signal \Lab_UT.scdp.q_RNIDHFGA_3\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_2\ : std_logic;
signal \Lab_UT.scdp.e2dData_2\ : std_logic;
signal \Lab_UT.scdp.N_59_i\ : std_logic;
signal \Lab_UT.scdp.pinst0.un12_pValidZ0Z_1\ : std_logic;
signal \Lab_UT.scdp.msBitsi.msBitsD_4\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_4\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_4_cascade_\ : std_logic;
signal \Lab_UT.scdp.q_RNIIAV0D_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.msBitsi.q_esr_RNI239EZ0Z_4\ : std_logic;
signal \ufifo.txdataDZ0Z_4\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_3\ : std_logic;
signal \Lab_UT.scdp.pValid_0\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_3_cascade_\ : std_logic;
signal \Lab_UT.scdp.lsBitsi.q_esr_RNI0TMAZ0Z_3\ : std_logic;
signal \Lab_UT.scdp.q_RNIRM8BD_3_cascade_\ : std_logic;
signal \ufifo.txdataDZ0Z_3\ : std_logic;
signal \Lab_UT.scdp.byteToDecrypt_0\ : std_logic;
signal \Lab_UT.scdp.byteToDecrypt_3\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_4\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_4\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_5\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_5\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_2\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_3\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_3\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_2\ : std_logic;
signal \ufifo.fifo.wraddrZ0Z_1\ : std_logic;
signal \ufifo.fifo.un1_emptyB_NE_0_cascade_\ : std_logic;
signal \ufifo.fifo.rdaddrZ0Z_1\ : std_logic;
signal \ufifo.tx_fsm.fifo_txdata_rdy\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \ufifo.fifo.un1_emptyB_NE_2\ : std_logic;
signal \ufifo.fifo.un1_emptyB_NE_1\ : std_logic;
signal \ufifo.fifo.un1_emptyB_NE_3\ : std_logic;
signal \ufifo.fifo.un1_emptyB_NE_4\ : std_logic;
signal \ufifo.emptyB_0_cascade_\ : std_logic;
signal \ufifo.tx_fsm.cstateZ0Z_1\ : std_logic;
signal \ufifo.tx_fsm.N_62_0_cascade_\ : std_logic;
signal \ufifo.popFifo\ : std_logic;
signal rst_i_3_i : std_logic;
signal \ufifo.emitcrlf_fsm.cstateZ0Z_0\ : std_logic;
signal \buart.Z_rx.bitcountlde_i_o2_0_cascade_\ : std_logic;
signal \buart.Z_rx.N_58_cascade_\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \buart.Z_rx.N_58\ : std_logic;
signal \buart.Z_rx.startbit_cascade_\ : std_logic;
signal \buart.Z_rx.ser_clk\ : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \buart.Z_rx.N_41_i_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \buart.Z_rx.N_45\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.N_43\ : std_logic;
signal \Lab_UT.dk.de_bigL_sxZ0\ : std_logic;
signal \Lab_UT.de_bigL_3\ : std_logic;
signal \Lab_UT.scctrl.g0_17_N_3LZ0Z3\ : std_logic;
signal \Lab_UT.de_bigL_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_17_N_2LZ0Z1\ : std_logic;
signal \Lab_UT.de_bigL_0\ : std_logic;
signal \buart__rx_bitcount_3\ : std_logic;
signal \buart__rx_bitcount_0\ : std_logic;
signal \buart__rx_bitcount_1\ : std_logic;
signal \buart__rx_bitcount_4\ : std_logic;
signal \buart.Z_rx.shifter_0_fast_RNI1CIH1Z0Z_2\ : std_logic;
signal \buart.Z_rx.bitcount_es_RNIF6D61Z0Z_4_cascade_\ : std_logic;
signal \Lab_UT_dk_de_bigD_0\ : std_logic;
signal \Lab_UT.dk.de_bigD_sxZ0\ : std_logic;
signal \Lab_UT_dk_de_bigD_0_cascade_\ : std_logic;
signal \Lab_UT.dk.de_bigD_1Z0Z_0\ : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_14\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_15\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_3\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_23\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28\ : std_logic;
signal \Lab_UT.scdp.prng_lfsr_7\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_5\ : std_logic;
signal \Lab_UT.scdp.d2eData_3_5_cascade_\ : std_logic;
signal \Lab_UT.scdp.e2dData_5\ : std_logic;
signal \Lab_UT.scdp.u0.byteToDecrypt_5\ : std_logic;
signal \Lab_UT.scdp.u0.byteToDecrypt_7\ : std_logic;
signal \Lab_UT.scdp.val_0_3\ : std_logic;
signal \Lab_UT.scdp.key1_7\ : std_logic;
signal \Lab_UT.scdp.key1_3\ : std_logic;
signal \ufifo.txDataValidDZ0\ : std_logic;
signal \ufifo.emitcrlf_fsm.cstate_srsts_sn_1\ : std_logic;
signal \ufifo.N_57_0_1_cascade_\ : std_logic;
signal \ufifo.tx_fsm.cstateZ0Z_4\ : std_logic;
signal \ufifo.tx_fsm.N_59_0\ : std_logic;
signal \buart__tx_uart_busy_0\ : std_logic;
signal \ufifo.emitcrlf_fsm.cstateZ0Z_1\ : std_logic;
signal \ufifo.emitcrlf_fsm.cstate_srsts_rn_0_1\ : std_logic;
signal \ufifo.tx_fsm.cstateZ0Z_5\ : std_logic;
signal \ufifo.crlfdone\ : std_logic;
signal \ufifo.tx_fsm.N_72_cascade_\ : std_logic;
signal \ufifo.cstate_0\ : std_logic;
signal \Lab_UT.dk.de_bigEZ0Z_2\ : std_logic;
signal \Lab_UT.scctrl.m24_e_4\ : std_logic;
signal \Lab_UT.dk.escKey_4_reti_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a7_1\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a3_2_cascade_\ : std_logic;
signal \Lab_UT.g0_i_a9_1_3_cascade_\ : std_logic;
signal \bu_rx_data_rdy_cascade_\ : std_logic;
signal \Lab_UT.scctrl.delay1\ : std_logic;
signal \Lab_UT.scctrl.delay2\ : std_logic;
signal \N_6\ : std_logic;
signal \Lab_UT.scdp.pinst1.un12_pValidZ0Z_1_cascade_\ : std_logic;
signal \Lab_UT.un7_pValid\ : std_logic;
signal \Lab_UT.un1_pValid\ : std_logic;
signal \Lab_UT.un7_pValid_cascade_\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_1_0_i_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_0_sqmuxa_4Z0Z_0\ : std_logic;
signal \Lab_UT.dk.de_bigEZ0Z_1\ : std_logic;
signal \Lab_UT_dk_de_bigD_6_cascade_\ : std_logic;
signal \Lab_UT.de_bigE_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_39_cascade_\ : std_logic;
signal \Lab_UT.scdp.a2b.N_50_cascade_\ : std_logic;
signal \Lab_UT.scdp.a2b.N_51\ : std_logic;
signal bu_rx_data_i_2_5 : std_logic;
signal \Lab_UT.scctrl.m24_e_5\ : std_logic;
signal \Lab_UT.scdp.a2b.N_50\ : std_logic;
signal bu_rx_data_3 : std_logic;
signal \Lab_UT.scdp.a2b.N_53_cascade_\ : std_logic;
signal \Lab_UT.scdp.N_39\ : std_logic;
signal \Lab_UT.scdp.byteToDecrypt_4\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_6\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsr_next_1_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_4\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_11\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_12\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_g\ : std_logic;
signal \Lab_UT.scdp.key3_0\ : std_logic;
signal \buart__rx_bitcount_2\ : std_logic;
signal \buart.Z_rx.bitcount_es_RNIGTPI1Z0Z_3\ : std_logic;
signal \Lab_UT.scdp.d2eData_0\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_0\ : std_logic;
signal \Lab_UT.scdp.lsBits_6\ : std_logic;
signal \Lab_UT.scdp.lsBitsD_4\ : std_logic;
signal \Lab_UT.scdp.N_48_i\ : std_logic;
signal \Lab_UT.scdp.N_52\ : std_logic;
signal \Lab_UT.scdp.msBitsD_3\ : std_logic;
signal \buart__tx_uart_busy_0_i\ : std_logic;
signal \buart.Z_tx.N_255\ : std_logic;
signal ufifo_utb_txdata_rdy_0 : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \Lab_UT.scctrl.delay3\ : std_logic;
signal \Lab_UT.scctrl.r4.delay4\ : std_logic;
signal \Lab_UT.scdp.u1.byteToDecrypt_2\ : std_logic;
signal \Lab_UT.scdp.key1_5\ : std_logic;
signal \Lab_UT.scdp.key1_1\ : std_logic;
signal \Lab_UT.scdp.key2_5\ : std_logic;
signal \Lab_UT.scdp.key3_5\ : std_logic;
signal \Lab_UT.scdp.key3_1\ : std_logic;
signal \Lab_UT.scdp.key1_0\ : std_logic;
signal \Lab_UT.scdp.key2_4\ : std_logic;
signal \Lab_UT.scdp.key3_4\ : std_logic;
signal \Lab_UT.sccEldByte\ : std_logic;
signal \Lab_UT.state_ret_6_RNIL97G01_0\ : std_logic;
signal \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_iZ0\ : std_logic;
signal \Lab_UT.scctrl.un1_state_inv_cascade_\ : std_logic;
signal \Lab_UT.scctrl.state_ret_12_RNIUQFKZ0_cascade_\ : std_logic;
signal \Lab_UT.state_ret_12_RNIMJCP8_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.delayload\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_1_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.un1_state_3_1_reti_cascade_\ : std_logic;
signal \Lab_UT.de_bigE_0\ : std_logic;
signal \Lab_UT.scctrl.g0_7_1_0\ : std_logic;
signal \Lab_UT.scctrl.g2_0_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_7_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1_0\ : std_logic;
signal \Lab_UT.scctrl.g2_2\ : std_logic;
signal \Lab_UT.scctrl.g1\ : std_logic;
signal \Lab_UT.sccDnibble1En\ : std_logic;
signal \Lab_UT.sccDnibble1En_cascade_\ : std_logic;
signal \Lab_UT.scdp.u0.sccDnibble1En_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_sqmuxa_3_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.state_retZ0Z_10\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_sqmuxa_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.nibbleInZ0Z1\ : std_logic;
signal \Lab_UT.scctrl.N_1_0_i\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_sqmuxa_3\ : std_logic;
signal \Lab_UT.scctrl.un6_sccDecrypt\ : std_logic;
signal \Lab_UT.de_bigE\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_i_a5_1_0\ : std_logic;
signal \Lab_UT.scctrl.EmsLoaded\ : std_logic;
signal \Lab_UT.scctrl.EmsLoaded_cascade_\ : std_logic;
signal \Lab_UT.sccElsBitsLd_cascade_\ : std_logic;
signal \Lab_UT.scdp.sccElsBitsLd_0\ : std_logic;
signal \Lab_UT.sccElsBitsLd\ : std_logic;
signal \Lab_UT.scdp.lsBitsi.lsBitsD_5\ : std_logic;
signal \Lab_UT_dk_de_cr_12_1_cascade_\ : std_logic;
signal \L4_PrintBuf_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_9_0\ : std_logic;
signal bu_rx_data_fast_0 : std_logic;
signal \buart__rx_shifter_0_fast_3\ : std_logic;
signal \Lab_UT.dk.un7_de_hex_xZ0Z0_cascade_\ : std_logic;
signal \Lab_UT.dk.un7_de_hex_0_cascade_\ : std_logic;
signal \Lab_UT.dk.un7_de_hex_0\ : std_logic;
signal \Lab_UT.un4_de_hex_cascade_\ : std_logic;
signal \buart__rx_shifter_0_fast_1\ : std_logic;
signal \buart__rx_shifter_ret_1_fast\ : std_logic;
signal \Lab_UT.scctrl.g0_i_o9_0Z0Z_2\ : std_logic;
signal \Lab_UT.dk.un4_de_hexZ0Z_1\ : std_logic;
signal bu_rx_data_i_3_4 : std_logic;
signal bu_rx_data_5 : std_logic;
signal bu_rx_data_4 : std_logic;
signal bu_rx_data_i_2_6 : std_logic;
signal \Lab_UT.un1_de_hex_2\ : std_logic;
signal \Lab_UT.un1_de_hex_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a9_3_4_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a9_3_5\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_0_a5_2_out_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_222_1\ : std_logic;
signal \Lab_UT.scctrl.next_state_3_sqmuxa_0\ : std_logic;
signal \Lab_UT.scdp.a2b.g1_1_a3_0Z0Z_0\ : std_logic;
signal \Lab_UT.scdp.key0_0\ : std_logic;
signal \Lab_UT.scdp.key0_2\ : std_logic;
signal \Lab_UT.scdp.key1_4\ : std_logic;
signal \Lab_UT.state_ret_13_RNIQ72741_0\ : std_logic;
signal \Lab_UT.scdp.key1_6\ : std_logic;
signal \Lab_UT.scctrl.next_state77_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_3_sqmuxa\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state77\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state77_2\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz_4\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz\ : std_logic;
signal \Lab_UT.scctrl.next_state76\ : std_logic;
signal \Lab_UT.scdp.key2_3\ : std_logic;
signal \Lab_UT.scdp.key2_6\ : std_logic;
signal \Lab_UT.state_ret_14_RNI416G41_0\ : std_logic;
signal \Lab_UT.scdp.key3_6\ : std_logic;
signal \Lab_UT.scdp.key3_2\ : std_logic;
signal \Lab_UT.state_2_RNI44QH41_0_2\ : std_logic;
signal \Lab_UT.scdp.key2_7\ : std_logic;
signal \Lab_UT.state_2_RNIF0RJ41_0_2\ : std_logic;
signal \Lab_UT.scdp.key3_3\ : std_logic;
signal \Lab_UT.state_ret_13_RNIHUNI41_0\ : std_logic;
signal \Lab_UT.state_ret_13_RNIHUNI41_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.key1_2\ : std_logic;
signal \Lab_UT.sccDecrypt_0\ : std_logic;
signal \Lab_UT.state_ret_12_RNIMJCP8_0\ : std_logic;
signal \Lab_UT.sccDnibble2En_cascade_\ : std_logic;
signal \resetGen_rst_0_iso\ : std_logic;
signal \Lab_UT.scdp.u1.sccDnibble2En_0\ : std_logic;
signal \Lab_UT.scdp.N_37\ : std_logic;
signal \Lab_UT.sccDnibble2En\ : std_logic;
signal \Lab_UT.scdp.byteToDecrypt_1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a9_0_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a9_1\ : std_logic;
signal \Lab_UT.scctrl.N_12_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_i_2\ : std_logic;
signal \Lab_UT.scctrl.G_23_0_a9_0_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a10_2_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.G_23_0_2\ : std_logic;
signal \Lab_UT.scctrl.N_2ctr\ : std_logic;
signal \Lab_UT.scctrl.g0_i_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_4\ : std_logic;
signal \Lab_UT.scctrl.N_10\ : std_logic;
signal \Lab_UT.scctrl.G_23_0_a9_4_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.G_23_0_3\ : std_logic;
signal \Lab_UT.scctrl.G_23_0_a9_3_1\ : std_logic;
signal \Lab_UT.scctrl.G_23_0_4\ : std_logic;
signal \Lab_UT.scctrl.G_23_0_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_3ctr\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a7_2_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_i_a5_4_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_8_0\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.state_i_3_fast_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_1_1_0\ : std_logic;
signal \Lab_UT.scdp.a2b.N_6_0\ : std_logic;
signal \Lab_UT.scctrl.g0_14_mb_rn_0\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_7_2\ : std_logic;
signal \Lab_UT.scctrl.state_i_3_fast_2\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_0_a5_0_0_3\ : std_logic;
signal \N_127_i_i_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_11_0\ : std_logic;
signal \Lab_UT.N_166_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_127_i_i_3\ : std_logic;
signal \Lab_UT.g1_i_a4_0_2_cascade_\ : std_logic;
signal \Lab_UT.next_state_3\ : std_logic;
signal \Lab_UT.g0_3_a3_0_4_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_8_0\ : std_logic;
signal \Lab_UT.scdp.a2b.g1_1_o2_0Z0Z_0\ : std_logic;
signal \Lab_UT.scdp.a2b.N_6_1_cascade_\ : std_logic;
signal \Lab_UT.scdp.a2b.g0_3_a3_0Z0Z_3\ : std_logic;
signal \Lab_UT.N_190\ : std_logic;
signal \Lab_UT.scctrl.N_6_3_0\ : std_logic;
signal \Lab_UT.scctrl.g0_1_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_2_0\ : std_logic;
signal \Lab_UT.scctrl.N_12_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_1_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_3_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.un6_sccDecrypt_0\ : std_logic;
signal \Lab_UT.scctrl.g1_1_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g2_0\ : std_logic;
signal \Lab_UT.scctrl.g0_1_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_1_3_1_cascade_\ : std_logic;
signal \Lab_UT.next_state_rst_1_3\ : std_logic;
signal \Lab_UT.next_state_rst_1_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_166_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_1_cascade_\ : std_logic;
signal led_c_2 : std_logic;
signal \Lab_UT.scctrl.g0_17_N_4LZ0Z5\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_3_N_6_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_i_2_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_2_0\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_3_N_6_1\ : std_logic;
signal \Lab_UT.g0_3_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a8_3_0\ : std_logic;
signal \Lab_UT.scctrl.N_6_3\ : std_logic;
signal \Lab_UT.scctrl.g0_i_1_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_0_1_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state75\ : std_logic;
signal \Lab_UT.scctrl.N_7_1\ : std_logic;
signal \Lab_UT.scctrl.N_223_2\ : std_logic;
signal \Lab_UT.scctrl.next_state73\ : std_logic;
signal \Lab_UT.scctrl.next_state73_cascade_\ : std_logic;
signal \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i\ : std_logic;
signal \Lab_UT.state_ret_3_RNII68F41_0_cascade_\ : std_logic;
signal \Lab_UT.scdp.key2_0\ : std_logic;
signal \Lab_UT.scdp.key2_1\ : std_logic;
signal \Lab_UT.state_ret_3_RNII68F41_0\ : std_logic;
signal \Lab_UT.scdp.key2_2\ : std_logic;
signal bu_rx_data_i_3_1 : std_logic;
signal \Lab_UT.scdp.key0_5\ : std_logic;
signal \Lab_UT.scdp.a2b.N_53\ : std_logic;
signal bu_rx_data_1 : std_logic;
signal bu_rx_data_2 : std_logic;
signal \Lab_UT.scdp.binValD_2\ : std_logic;
signal \Lab_UT.scdp.key0_6\ : std_logic;
signal \Lab_UT.scdp.binValD_0\ : std_logic;
signal \Lab_UT.scdp.key0_4\ : std_logic;
signal \Lab_UT.state_ret_RNIUV0941_0\ : std_logic;
signal \Lab_UT.scdp.key0_7\ : std_logic;
signal \Lab_UT.scdp.binValD_1\ : std_logic;
signal \Lab_UT.scdp.key0_1\ : std_logic;
signal \Lab_UT.scdp.binValD_3\ : std_logic;
signal \Lab_UT.scdp.binVal_ValidD\ : std_logic;
signal \Lab_UT.state_0_RNIKFK051_0_1\ : std_logic;
signal \Lab_UT.scdp.key0_3\ : std_logic;
signal \Lab_UT.scctrl.next_state74\ : std_logic;
signal \G_23_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_12_1\ : std_logic;
signal \Lab_UT.scctrl.N_5_0\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_a8_3_1_0\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_a8_2_1_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_3_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_13\ : std_logic;
signal \Lab_UT.scctrl.g0_i_1\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_2\ : std_logic;
signal \Lab_UT.scctrl.g0_16_mb_sn\ : std_logic;
signal \Lab_UT.scctrl.g0_16_mb_rn_0\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_3_0\ : std_logic;
signal \Lab_UT_dk_de_cr_12_1\ : std_logic;
signal \ufifo.emptyB_0\ : std_logic;
signal bu_rx_data_0 : std_logic;
signal \ufifo.tx_fsm.N_60_0\ : std_logic;
signal \Lab_UT.scctrl.N_127_i_i_a6_0_0\ : std_logic;
signal \Lab_UT.scctrl.N_11\ : std_logic;
signal \Lab_UT.scctrl.G_21_i_a7_1_1\ : std_logic;
signal \Lab_UT.m61_i_a2_2\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_0_0\ : std_logic;
signal \Lab_UT.N_5_cascade_\ : std_logic;
signal \Lab_UT.g0_i_5\ : std_logic;
signal \Lab_UT.scctrl.g0_14_mb_sn\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_1_1\ : std_logic;
signal \Lab_UT.scctrl.N_14\ : std_logic;
signal \Lab_UT.scdp.a2b.g0_iZ0Z_4\ : std_logic;
signal \Lab_UT.N_5\ : std_logic;
signal \Lab_UT.scdp.a2b.g0_iZ0Z_8_cascade_\ : std_logic;
signal \Lab_UT.scdp.a2b.g0_3_a3_6\ : std_logic;
signal \Lab_UT.de_cr_2\ : std_logic;
signal \Lab_UT.de_cr_6_0\ : std_logic;
signal \Lab_UT.g0_i_a5_1_3_cascade_\ : std_logic;
signal \Lab_UT.scdp.a2b.N_9_1\ : std_logic;
signal \Lab_UT.scdp.a2b.g1_1_0_1\ : std_logic;
signal \Lab_UT.scctrl.g0_1_3_1\ : std_logic;
signal \Lab_UT.scctrl.N_127_i_i_o6_0_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_127_i_i_a6_1\ : std_logic;
signal \Lab_UT.scctrl.N_190_0_0\ : std_logic;
signal \Lab_UT.next_state_rst_0_5\ : std_logic;
signal \Lab_UT.scdp.a2b.N_6_4\ : std_logic;
signal \Lab_UT.state_ret_8_rep1_RNIHA8U3\ : std_logic;
signal \Lab_UT.N_182\ : std_logic;
signal \Lab_UT.scdp.a2b.g0_iZ0Z_9\ : std_logic;
signal \Lab_UT.state_2_RNI3PVB9_2\ : std_logic;
signal \Lab_UT.scctrl.N_182_0\ : std_logic;
signal \Lab_UT.scctrl.N_166_0_1\ : std_logic;
signal bu_rx_data_0_rep1 : std_logic;
signal \Lab_UT.scctrl.next_state_1_i_o2_0_d_1_cascade_\ : std_logic;
signal \buart__rx_shifter_0_fast_2\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_3_N_5L8Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT_dk_de_bigD_6\ : std_logic;
signal \shifter_0_fast_RNI639J4_2\ : std_logic;
signal \Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433_cascade_\ : std_logic;
signal \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0\ : std_logic;
signal \Lab_UT.de_bigD\ : std_logic;
signal \Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433\ : std_logic;
signal \Lab_UT.de_bigL\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_i_o2_0_d_1\ : std_logic;
signal \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0Z_2\ : std_logic;
signal bu_rx_data_6 : std_logic;
signal bu_rx_data_7 : std_logic;
signal \resetGen_escKey_4\ : std_logic;
signal \N_41_i_g\ : std_logic;
signal \Lab_UT.scctrl.g0_2_1\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_3_N_6_0\ : std_logic;
signal \Lab_UT.scctrl.g1_0_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_1_3\ : std_logic;
signal \Lab_UT.scctrl.g0_1_0_0\ : std_logic;
signal rst_i_3_rep2 : std_logic;
signal \Lab_UT.state_ret_8_rep1_RNIJDTUE_1\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_0_5_0_cascade_\ : std_logic;
signal \Lab_UT.scctrl.stateZ0Z_3\ : std_logic;
signal rst_i_3_rep1 : std_logic;
signal \Lab_UT.scctrl.g0_i_a8_1\ : std_logic;
signal \Lab_UT.scctrl.g0_i_0_0\ : std_logic;
signal \Lab_UT.scctrl.g0_7_3\ : std_logic;
signal \Lab_UT.scctrl.g0_7_2\ : std_logic;
signal \Lab_UT.scctrl.g2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1_1\ : std_logic;
signal \Lab_UT.scctrl.g0_1_0\ : std_logic;
signal \Lab_UT.scctrl.N_222i_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_223_1_reti\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_2\ : std_logic;
signal \Lab_UT.scctrl.N_223_2_reti\ : std_logic;
signal \Lab_UT.next_state_rst_2_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_3\ : std_logic;
signal \Lab_UT.scctrl.N_8\ : std_logic;
signal \Lab_UT.scctrl.g0_i_4_0_cascade_\ : std_logic;
signal led_c_0 : std_logic;
signal \Lab_UT.scctrl.N_8_1\ : std_logic;
signal \Lab_UT.scctrl.N_8_3\ : std_logic;
signal \Lab_UT.scctrl.g0_18_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_stateZ0Z_2\ : std_logic;
signal \Lab_UT.scctrl.next_stateZ0Z_2_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_6_2\ : std_logic;
signal \Lab_UT.scctrl.g0_i_3_1\ : std_logic;
signal next_state_1 : std_logic;
signal \Lab_UT.scctrl.g0_i_m4_1_1\ : std_logic;
signal \Lab_UT.scctrl.N_9\ : std_logic;
signal \Lab_UT.scctrl.g1_i_a7_1\ : std_logic;
signal \Lab_UT.scctrl.next_state_0_3\ : std_logic;
signal \Lab_UT.scctrl.next_state_1_0_3\ : std_logic;
signal \Lab_UT.scctrl.next_state_i_3_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_state71\ : std_logic;
signal \Lab_UT.scctrl.next_state72\ : std_logic;
signal \Lab_UT.scctrl.g4_1\ : std_logic;
signal \Lab_UT.sccEmsBitsSl\ : std_logic;
signal \Lab_UT.scctrl.g2\ : std_logic;
signal \Lab_UT.scctrl.next_state_rst_3\ : std_logic;
signal \resetGen_rst_0_iso_g\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_a8_0_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_20\ : std_logic;
signal \Lab_UT.scctrl.G_38_0_a3_0_4_cascade_\ : std_logic;
signal \Lab_UT.scctrl.next_stateZ0Z_0\ : std_logic;
signal \Lab_UT.scctrl.G_38_0_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_7_0\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_0\ : std_logic;
signal \Lab_UT.scdp.a2b.g0_i_a9_1\ : std_logic;
signal \Lab_UT.scdp.a2b.g0_iZ0Z_1_cascade_\ : std_logic;
signal \Lab_UT.scdp.a2b.g0_iZ0Z_2\ : std_logic;
signal \Lab_UT.scctrl.g0_7_a13_1_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_7_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g0_6\ : std_logic;
signal rst : std_logic;
signal \Lab_UT.scctrl.g1_i_a7_2Z0Z_3\ : std_logic;
signal \Lab_UT.scctrl.N_10_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.g1_i_2\ : std_logic;
signal \Lab_UT.scctrl.N_7_4\ : std_logic;
signal \Lab_UT.un1_de_hex\ : std_logic;
signal \Lab_UT.scctrl.G_21_i_a7_0\ : std_logic;
signal \Lab_UT.un4_de_hex\ : std_logic;
signal \Lab_UT.scctrl.N_11_1\ : std_logic;
signal \Lab_UT.scctrl.N_12_2\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_a4_1_cascade_\ : std_logic;
signal \Lab_UT.scctrl.G_21_i_a7_0_1\ : std_logic;
signal \Lab_UT.scctrl.N_9_2\ : std_logic;
signal \Lab_UT.scctrl.G_21_i_2\ : std_logic;
signal \Lab_UT.scctrl.N_8_2\ : std_logic;
signal \Lab_UT.state_i_3_0_rep1\ : std_logic;
signal \Lab_UT.state_i_3_2_rep1\ : std_logic;
signal \Lab_UT.scctrl.g0_1_4_1\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a7_0_1_cascade_\ : std_logic;
signal \Lab_UT.de_hex_0\ : std_logic;
signal \Lab_UT.scctrl.N_10_0\ : std_logic;
signal \Lab_UT.un1_state_3_1\ : std_logic;
signal \L4_PrintBuf\ : std_logic;
signal \Lab_UT.scctrl.m26_i_o4_1_2\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_o3_0_0_cascade_\ : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \Lab_UT.scctrl.N_6_5_cascade_\ : std_logic;
signal \Lab_UT.scctrl.N_5_2\ : std_logic;
signal \Lab_UT.scctrl.N_8_4\ : std_logic;
signal \Lab_UT.scctrl.N_4ctr\ : std_logic;
signal \Lab_UT.scctrl.G_23_0_a9_1\ : std_logic;
signal \Lab_UT.state_i_3_1\ : std_logic;
signal \Lab_UT.scctrl.g0_i_a8_4_1\ : std_logic;
signal \Lab_UT.scctrl.next_state_0_2\ : std_logic;
signal rst_i_3 : std_logic;
signal \Lab_UT_scctrl_N_221_0\ : std_logic;
signal \Lab_UT.scctrl.G_21_i_0\ : std_logic;
signal \Lab_UT.state_i_3_2\ : std_logic;
signal \Lab_UT.state_2\ : std_logic;
signal \Lab_UT.state_0\ : std_logic;
signal \Lab_UT.scctrl.g0_i_7_1\ : std_logic;
signal rst_i_3_reti : std_logic;
signal clk_g : std_logic;
signal \Lab_UT.scctrl.g2_1\ : std_logic;
signal \Lab_UT.state_i_3_2_rep2\ : std_logic;
signal \Lab_UT.state_i_3_3\ : std_logic;
signal \Lab_UT.scctrl.state_i_3_0_rep2\ : std_logic;
signal rst_i_3_fast : std_logic;
signal \Lab_UT.scctrl.g1_i_0\ : std_logic;
signal \Lab_UT.state_i_3_0\ : std_logic;
signal \Lab_UT.scctrl.g0_0_i_a8_3_1\ : std_logic;
signal \Lab_UT.state_1\ : std_logic;
signal \Lab_UT.scctrl.state_1_RNO_3Z0Z_0\ : std_logic;
signal \Lab_UT.scctrl.N_13_0\ : std_logic;
signal \Lab_UT.N_191\ : std_logic;
signal \Lab_UT.scctrl.G_24_i_a4_0_1\ : std_logic;
signal \Lab_UT.next_state_1_0_0_3\ : std_logic;
signal \Lab_UT.scctrl.N_10_2\ : std_logic;
signal \Lab_UT.N_169_0\ : std_logic;
signal \Lab_UT.scctrl.N_223_1\ : std_logic;
signal led_c_4 : std_logic;
signal \_gnd_net_\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \ufifo.fifo.sb_ram512x8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \ufifo.fifo.sb_ram512x8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \ufifo.fifo.sb_ram512x8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \ufifo.fifo.sb_ram512x8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    led <= led_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    \ufifo.fifo.fifo_txdata_7\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(14);
    \ufifo.fifo.fifo_txdata_6\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(12);
    \ufifo.fifo.fifo_txdata_5\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(10);
    \ufifo.fifo.fifo_txdata_4\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(8);
    \ufifo.fifo.fifo_txdata_3\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(6);
    \ufifo.fifo.fifo_txdata_2\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(4);
    \ufifo.fifo.fifo_txdata_1\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(2);
    \ufifo.fifo.fifo_txdata_0\ <= \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\(0);
    \ufifo.fifo.sb_ram512x8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__8587\&\N__8704\&\N__8644\&\N__9721\&\N__9781\&\N__9664\&\N__9604\&\N__9544\&\N__8527\;
    \ufifo.fifo.sb_ram512x8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__8560\&\N__8674\&\N__8734\&\N__9751\&\N__9808\&\N__9634\&\N__9691\&\N__9574\&\N__8614\;
    \ufifo.fifo.sb_ram512x8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \ufifo.fifo.sb_ram512x8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__8827\&'0'&\N__8983\&'0'&\N__9415\&'0'&\N__9868\&'0'&\N__9193\&'0'&\N__9010\&'0'&\N__8833\;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \ufifo.fifo.sb_ram512x8_inst_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \ufifo.fifo.sb_ram512x8_inst_physical_RDATA_wire\,
            RADDR => \ufifo.fifo.sb_ram512x8_inst_physical_RADDR_wire\,
            WADDR => \ufifo.fifo.sb_ram512x8_inst_physical_WADDR_wire\,
            MASK => \ufifo.fifo.sb_ram512x8_inst_physical_MASK_wire\,
            WDATA => \ufifo.fifo.sb_ram512x8_inst_physical_WDATA_wire\,
            RCLKE => \N__10025\,
            RCLK => \N__22671\,
            RE => \N__10026\,
            WCLKE => \N__11091\,
            WCLK => \N__22670\,
            WE => \N__11092\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \latticehx1k_pll_inst.clk\,
            REFERENCECLK => \N__7825\,
            RESETB => \N__13966\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23195\,
            DIN => \N__23194\,
            DOUT => \N__23193\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23195\,
            PADOUT => \N__23194\,
            PADIN => \N__23193\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21214\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23186\,
            DIN => \N__23185\,
            DOUT => \N__23184\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23186\,
            PADOUT => \N__23185\,
            PADIN => \N__23184\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17807\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23177\,
            DIN => \N__23176\,
            DOUT => \N__23175\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23177\,
            PADOUT => \N__23176\,
            PADIN => \N__23175\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23168\,
            DIN => \N__23167\,
            DOUT => \N__23166\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23168\,
            PADOUT => \N__23167\,
            PADIN => \N__23166\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17808\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23159\,
            DIN => \N__23158\,
            DOUT => \N__23157\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23159\,
            PADOUT => \N__23158\,
            PADIN => \N__23157\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__22662\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23150\,
            DIN => \N__23149\,
            DOUT => \N__23148\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__23150\,
            PADOUT => \N__23149\,
            PADIN => \N__23148\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23141\,
            DIN => \N__23140\,
            DOUT => \N__23139\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23141\,
            PADOUT => \N__23140\,
            PADIN => \N__23139\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23132\,
            DIN => \N__23131\,
            DOUT => \N__23130\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23132\,
            PADOUT => \N__23131\,
            PADIN => \N__23130\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8107\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23123\,
            DIN => \N__23122\,
            DOUT => \N__23121\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23123\,
            PADOUT => \N__23122\,
            PADIN => \N__23121\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23114\,
            DIN => \N__23113\,
            DOUT => \N__23112\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23114\,
            PADOUT => \N__23113\,
            PADIN => \N__23112\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14672\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__23095\,
            I => \N__23083\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__23094\,
            I => \N__23080\
        );

    \I__5741\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23069\
        );

    \I__5740\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23066\
        );

    \I__5739\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23057\
        );

    \I__5738\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23057\
        );

    \I__5737\ : CascadeMux
    port map (
            O => \N__23089\,
            I => \N__23054\
        );

    \I__5736\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23048\
        );

    \I__5735\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23045\
        );

    \I__5734\ : InMux
    port map (
            O => \N__23086\,
            I => \N__23042\
        );

    \I__5733\ : InMux
    port map (
            O => \N__23083\,
            I => \N__23039\
        );

    \I__5732\ : InMux
    port map (
            O => \N__23080\,
            I => \N__23036\
        );

    \I__5731\ : InMux
    port map (
            O => \N__23079\,
            I => \N__23031\
        );

    \I__5730\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23031\
        );

    \I__5729\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23026\
        );

    \I__5728\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23026\
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__23075\,
            I => \N__23023\
        );

    \I__5726\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23015\
        );

    \I__5725\ : CascadeMux
    port map (
            O => \N__23073\,
            I => \N__23012\
        );

    \I__5724\ : CascadeMux
    port map (
            O => \N__23072\,
            I => \N__23008\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__23069\,
            I => \N__23003\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__23066\,
            I => \N__23003\
        );

    \I__5721\ : InMux
    port map (
            O => \N__23065\,
            I => \N__22998\
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__23064\,
            I => \N__22995\
        );

    \I__5719\ : InMux
    port map (
            O => \N__23063\,
            I => \N__22988\
        );

    \I__5718\ : InMux
    port map (
            O => \N__23062\,
            I => \N__22988\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__23057\,
            I => \N__22985\
        );

    \I__5716\ : InMux
    port map (
            O => \N__23054\,
            I => \N__22976\
        );

    \I__5715\ : InMux
    port map (
            O => \N__23053\,
            I => \N__22976\
        );

    \I__5714\ : InMux
    port map (
            O => \N__23052\,
            I => \N__22976\
        );

    \I__5713\ : InMux
    port map (
            O => \N__23051\,
            I => \N__22976\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__23048\,
            I => \N__22971\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__23045\,
            I => \N__22971\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__23042\,
            I => \N__22968\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__23039\,
            I => \N__22961\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__23036\,
            I => \N__22961\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__23031\,
            I => \N__22961\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__23026\,
            I => \N__22958\
        );

    \I__5705\ : InMux
    port map (
            O => \N__23023\,
            I => \N__22950\
        );

    \I__5704\ : InMux
    port map (
            O => \N__23022\,
            I => \N__22950\
        );

    \I__5703\ : InMux
    port map (
            O => \N__23021\,
            I => \N__22947\
        );

    \I__5702\ : InMux
    port map (
            O => \N__23020\,
            I => \N__22944\
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__23019\,
            I => \N__22941\
        );

    \I__5700\ : InMux
    port map (
            O => \N__23018\,
            I => \N__22938\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__23015\,
            I => \N__22935\
        );

    \I__5698\ : InMux
    port map (
            O => \N__23012\,
            I => \N__22932\
        );

    \I__5697\ : InMux
    port map (
            O => \N__23011\,
            I => \N__22927\
        );

    \I__5696\ : InMux
    port map (
            O => \N__23008\,
            I => \N__22927\
        );

    \I__5695\ : IoSpan4Mux
    port map (
            O => \N__23003\,
            I => \N__22924\
        );

    \I__5694\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22921\
        );

    \I__5693\ : InMux
    port map (
            O => \N__23001\,
            I => \N__22916\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__22998\,
            I => \N__22913\
        );

    \I__5691\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22910\
        );

    \I__5690\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22907\
        );

    \I__5689\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22904\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__22988\,
            I => \N__22891\
        );

    \I__5687\ : Span4Mux_h
    port map (
            O => \N__22985\,
            I => \N__22891\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__22976\,
            I => \N__22891\
        );

    \I__5685\ : Span4Mux_v
    port map (
            O => \N__22971\,
            I => \N__22891\
        );

    \I__5684\ : Span4Mux_v
    port map (
            O => \N__22968\,
            I => \N__22891\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__22961\,
            I => \N__22891\
        );

    \I__5682\ : Span4Mux_h
    port map (
            O => \N__22958\,
            I => \N__22888\
        );

    \I__5681\ : InMux
    port map (
            O => \N__22957\,
            I => \N__22881\
        );

    \I__5680\ : InMux
    port map (
            O => \N__22956\,
            I => \N__22881\
        );

    \I__5679\ : InMux
    port map (
            O => \N__22955\,
            I => \N__22881\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22874\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__22947\,
            I => \N__22874\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__22944\,
            I => \N__22874\
        );

    \I__5675\ : InMux
    port map (
            O => \N__22941\,
            I => \N__22871\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__22938\,
            I => \N__22866\
        );

    \I__5673\ : Span4Mux_h
    port map (
            O => \N__22935\,
            I => \N__22866\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__22932\,
            I => \N__22863\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__22927\,
            I => \N__22860\
        );

    \I__5670\ : IoSpan4Mux
    port map (
            O => \N__22924\,
            I => \N__22857\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__22921\,
            I => \N__22854\
        );

    \I__5668\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22849\
        );

    \I__5667\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22849\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22846\
        );

    \I__5665\ : Span4Mux_v
    port map (
            O => \N__22913\,
            I => \N__22835\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__22910\,
            I => \N__22835\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__22907\,
            I => \N__22835\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__22904\,
            I => \N__22835\
        );

    \I__5661\ : Span4Mux_v
    port map (
            O => \N__22891\,
            I => \N__22835\
        );

    \I__5660\ : Span4Mux_v
    port map (
            O => \N__22888\,
            I => \N__22828\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__22881\,
            I => \N__22828\
        );

    \I__5658\ : Span4Mux_h
    port map (
            O => \N__22874\,
            I => \N__22828\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__22871\,
            I => \N__22817\
        );

    \I__5656\ : Span4Mux_v
    port map (
            O => \N__22866\,
            I => \N__22817\
        );

    \I__5655\ : Span4Mux_h
    port map (
            O => \N__22863\,
            I => \N__22817\
        );

    \I__5654\ : Span4Mux_h
    port map (
            O => \N__22860\,
            I => \N__22817\
        );

    \I__5653\ : Span4Mux_s1_h
    port map (
            O => \N__22857\,
            I => \N__22817\
        );

    \I__5652\ : Span12Mux_s1_h
    port map (
            O => \N__22854\,
            I => \N__22814\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__22849\,
            I => \Lab_UT.state_0\
        );

    \I__5650\ : Odrv12
    port map (
            O => \N__22846\,
            I => \Lab_UT.state_0\
        );

    \I__5649\ : Odrv4
    port map (
            O => \N__22835\,
            I => \Lab_UT.state_0\
        );

    \I__5648\ : Odrv4
    port map (
            O => \N__22828\,
            I => \Lab_UT.state_0\
        );

    \I__5647\ : Odrv4
    port map (
            O => \N__22817\,
            I => \Lab_UT.state_0\
        );

    \I__5646\ : Odrv12
    port map (
            O => \N__22814\,
            I => \Lab_UT.state_0\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__22801\,
            I => \N__22798\
        );

    \I__5644\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22795\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__22795\,
            I => \N__22792\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__22792\,
            I => \Lab_UT.scctrl.g0_i_7_1\
        );

    \I__5641\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22785\
        );

    \I__5640\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22782\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__22785\,
            I => \N__22775\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__22782\,
            I => \N__22775\
        );

    \I__5637\ : InMux
    port map (
            O => \N__22781\,
            I => \N__22772\
        );

    \I__5636\ : InMux
    port map (
            O => \N__22780\,
            I => \N__22769\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__22775\,
            I => \N__22758\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__22772\,
            I => \N__22753\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__22769\,
            I => \N__22753\
        );

    \I__5632\ : InMux
    port map (
            O => \N__22768\,
            I => \N__22748\
        );

    \I__5631\ : InMux
    port map (
            O => \N__22767\,
            I => \N__22748\
        );

    \I__5630\ : CascadeMux
    port map (
            O => \N__22766\,
            I => \N__22745\
        );

    \I__5629\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22737\
        );

    \I__5628\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22737\
        );

    \I__5627\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22737\
        );

    \I__5626\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22734\
        );

    \I__5625\ : InMux
    port map (
            O => \N__22761\,
            I => \N__22731\
        );

    \I__5624\ : Span4Mux_h
    port map (
            O => \N__22758\,
            I => \N__22724\
        );

    \I__5623\ : Span4Mux_v
    port map (
            O => \N__22753\,
            I => \N__22724\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__22748\,
            I => \N__22724\
        );

    \I__5621\ : InMux
    port map (
            O => \N__22745\,
            I => \N__22719\
        );

    \I__5620\ : InMux
    port map (
            O => \N__22744\,
            I => \N__22719\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__22737\,
            I => \N__22716\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__22734\,
            I => \N__22711\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__22731\,
            I => \N__22711\
        );

    \I__5616\ : Span4Mux_h
    port map (
            O => \N__22724\,
            I => \N__22708\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__22719\,
            I => rst_i_3_reti
        );

    \I__5614\ : Odrv12
    port map (
            O => \N__22716\,
            I => rst_i_3_reti
        );

    \I__5613\ : Odrv12
    port map (
            O => \N__22711\,
            I => rst_i_3_reti
        );

    \I__5612\ : Odrv4
    port map (
            O => \N__22708\,
            I => rst_i_3_reti
        );

    \I__5611\ : ClkMux
    port map (
            O => \N__22699\,
            I => \N__22441\
        );

    \I__5610\ : ClkMux
    port map (
            O => \N__22698\,
            I => \N__22441\
        );

    \I__5609\ : ClkMux
    port map (
            O => \N__22697\,
            I => \N__22441\
        );

    \I__5608\ : ClkMux
    port map (
            O => \N__22696\,
            I => \N__22441\
        );

    \I__5607\ : ClkMux
    port map (
            O => \N__22695\,
            I => \N__22441\
        );

    \I__5606\ : ClkMux
    port map (
            O => \N__22694\,
            I => \N__22441\
        );

    \I__5605\ : ClkMux
    port map (
            O => \N__22693\,
            I => \N__22441\
        );

    \I__5604\ : ClkMux
    port map (
            O => \N__22692\,
            I => \N__22441\
        );

    \I__5603\ : ClkMux
    port map (
            O => \N__22691\,
            I => \N__22441\
        );

    \I__5602\ : ClkMux
    port map (
            O => \N__22690\,
            I => \N__22441\
        );

    \I__5601\ : ClkMux
    port map (
            O => \N__22689\,
            I => \N__22441\
        );

    \I__5600\ : ClkMux
    port map (
            O => \N__22688\,
            I => \N__22441\
        );

    \I__5599\ : ClkMux
    port map (
            O => \N__22687\,
            I => \N__22441\
        );

    \I__5598\ : ClkMux
    port map (
            O => \N__22686\,
            I => \N__22441\
        );

    \I__5597\ : ClkMux
    port map (
            O => \N__22685\,
            I => \N__22441\
        );

    \I__5596\ : ClkMux
    port map (
            O => \N__22684\,
            I => \N__22441\
        );

    \I__5595\ : ClkMux
    port map (
            O => \N__22683\,
            I => \N__22441\
        );

    \I__5594\ : ClkMux
    port map (
            O => \N__22682\,
            I => \N__22441\
        );

    \I__5593\ : ClkMux
    port map (
            O => \N__22681\,
            I => \N__22441\
        );

    \I__5592\ : ClkMux
    port map (
            O => \N__22680\,
            I => \N__22441\
        );

    \I__5591\ : ClkMux
    port map (
            O => \N__22679\,
            I => \N__22441\
        );

    \I__5590\ : ClkMux
    port map (
            O => \N__22678\,
            I => \N__22441\
        );

    \I__5589\ : ClkMux
    port map (
            O => \N__22677\,
            I => \N__22441\
        );

    \I__5588\ : ClkMux
    port map (
            O => \N__22676\,
            I => \N__22441\
        );

    \I__5587\ : ClkMux
    port map (
            O => \N__22675\,
            I => \N__22441\
        );

    \I__5586\ : ClkMux
    port map (
            O => \N__22674\,
            I => \N__22441\
        );

    \I__5585\ : ClkMux
    port map (
            O => \N__22673\,
            I => \N__22441\
        );

    \I__5584\ : ClkMux
    port map (
            O => \N__22672\,
            I => \N__22441\
        );

    \I__5583\ : ClkMux
    port map (
            O => \N__22671\,
            I => \N__22441\
        );

    \I__5582\ : ClkMux
    port map (
            O => \N__22670\,
            I => \N__22441\
        );

    \I__5581\ : ClkMux
    port map (
            O => \N__22669\,
            I => \N__22441\
        );

    \I__5580\ : ClkMux
    port map (
            O => \N__22668\,
            I => \N__22441\
        );

    \I__5579\ : ClkMux
    port map (
            O => \N__22667\,
            I => \N__22441\
        );

    \I__5578\ : ClkMux
    port map (
            O => \N__22666\,
            I => \N__22441\
        );

    \I__5577\ : ClkMux
    port map (
            O => \N__22665\,
            I => \N__22441\
        );

    \I__5576\ : ClkMux
    port map (
            O => \N__22664\,
            I => \N__22441\
        );

    \I__5575\ : ClkMux
    port map (
            O => \N__22663\,
            I => \N__22441\
        );

    \I__5574\ : ClkMux
    port map (
            O => \N__22662\,
            I => \N__22441\
        );

    \I__5573\ : ClkMux
    port map (
            O => \N__22661\,
            I => \N__22441\
        );

    \I__5572\ : ClkMux
    port map (
            O => \N__22660\,
            I => \N__22441\
        );

    \I__5571\ : ClkMux
    port map (
            O => \N__22659\,
            I => \N__22441\
        );

    \I__5570\ : ClkMux
    port map (
            O => \N__22658\,
            I => \N__22441\
        );

    \I__5569\ : ClkMux
    port map (
            O => \N__22657\,
            I => \N__22441\
        );

    \I__5568\ : ClkMux
    port map (
            O => \N__22656\,
            I => \N__22441\
        );

    \I__5567\ : ClkMux
    port map (
            O => \N__22655\,
            I => \N__22441\
        );

    \I__5566\ : ClkMux
    port map (
            O => \N__22654\,
            I => \N__22441\
        );

    \I__5565\ : ClkMux
    port map (
            O => \N__22653\,
            I => \N__22441\
        );

    \I__5564\ : ClkMux
    port map (
            O => \N__22652\,
            I => \N__22441\
        );

    \I__5563\ : ClkMux
    port map (
            O => \N__22651\,
            I => \N__22441\
        );

    \I__5562\ : ClkMux
    port map (
            O => \N__22650\,
            I => \N__22441\
        );

    \I__5561\ : ClkMux
    port map (
            O => \N__22649\,
            I => \N__22441\
        );

    \I__5560\ : ClkMux
    port map (
            O => \N__22648\,
            I => \N__22441\
        );

    \I__5559\ : ClkMux
    port map (
            O => \N__22647\,
            I => \N__22441\
        );

    \I__5558\ : ClkMux
    port map (
            O => \N__22646\,
            I => \N__22441\
        );

    \I__5557\ : ClkMux
    port map (
            O => \N__22645\,
            I => \N__22441\
        );

    \I__5556\ : ClkMux
    port map (
            O => \N__22644\,
            I => \N__22441\
        );

    \I__5555\ : ClkMux
    port map (
            O => \N__22643\,
            I => \N__22441\
        );

    \I__5554\ : ClkMux
    port map (
            O => \N__22642\,
            I => \N__22441\
        );

    \I__5553\ : ClkMux
    port map (
            O => \N__22641\,
            I => \N__22441\
        );

    \I__5552\ : ClkMux
    port map (
            O => \N__22640\,
            I => \N__22441\
        );

    \I__5551\ : ClkMux
    port map (
            O => \N__22639\,
            I => \N__22441\
        );

    \I__5550\ : ClkMux
    port map (
            O => \N__22638\,
            I => \N__22441\
        );

    \I__5549\ : ClkMux
    port map (
            O => \N__22637\,
            I => \N__22441\
        );

    \I__5548\ : ClkMux
    port map (
            O => \N__22636\,
            I => \N__22441\
        );

    \I__5547\ : ClkMux
    port map (
            O => \N__22635\,
            I => \N__22441\
        );

    \I__5546\ : ClkMux
    port map (
            O => \N__22634\,
            I => \N__22441\
        );

    \I__5545\ : ClkMux
    port map (
            O => \N__22633\,
            I => \N__22441\
        );

    \I__5544\ : ClkMux
    port map (
            O => \N__22632\,
            I => \N__22441\
        );

    \I__5543\ : ClkMux
    port map (
            O => \N__22631\,
            I => \N__22441\
        );

    \I__5542\ : ClkMux
    port map (
            O => \N__22630\,
            I => \N__22441\
        );

    \I__5541\ : ClkMux
    port map (
            O => \N__22629\,
            I => \N__22441\
        );

    \I__5540\ : ClkMux
    port map (
            O => \N__22628\,
            I => \N__22441\
        );

    \I__5539\ : ClkMux
    port map (
            O => \N__22627\,
            I => \N__22441\
        );

    \I__5538\ : ClkMux
    port map (
            O => \N__22626\,
            I => \N__22441\
        );

    \I__5537\ : ClkMux
    port map (
            O => \N__22625\,
            I => \N__22441\
        );

    \I__5536\ : ClkMux
    port map (
            O => \N__22624\,
            I => \N__22441\
        );

    \I__5535\ : ClkMux
    port map (
            O => \N__22623\,
            I => \N__22441\
        );

    \I__5534\ : ClkMux
    port map (
            O => \N__22622\,
            I => \N__22441\
        );

    \I__5533\ : ClkMux
    port map (
            O => \N__22621\,
            I => \N__22441\
        );

    \I__5532\ : ClkMux
    port map (
            O => \N__22620\,
            I => \N__22441\
        );

    \I__5531\ : ClkMux
    port map (
            O => \N__22619\,
            I => \N__22441\
        );

    \I__5530\ : ClkMux
    port map (
            O => \N__22618\,
            I => \N__22441\
        );

    \I__5529\ : ClkMux
    port map (
            O => \N__22617\,
            I => \N__22441\
        );

    \I__5528\ : ClkMux
    port map (
            O => \N__22616\,
            I => \N__22441\
        );

    \I__5527\ : ClkMux
    port map (
            O => \N__22615\,
            I => \N__22441\
        );

    \I__5526\ : ClkMux
    port map (
            O => \N__22614\,
            I => \N__22441\
        );

    \I__5525\ : GlobalMux
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__5524\ : gio2CtrlBuf
    port map (
            O => \N__22438\,
            I => clk_g
        );

    \I__5523\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22432\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__5521\ : Span4Mux_h
    port map (
            O => \N__22429\,
            I => \N__22426\
        );

    \I__5520\ : Odrv4
    port map (
            O => \N__22426\,
            I => \Lab_UT.scctrl.g2_1\
        );

    \I__5519\ : InMux
    port map (
            O => \N__22423\,
            I => \N__22417\
        );

    \I__5518\ : CascadeMux
    port map (
            O => \N__22422\,
            I => \N__22411\
        );

    \I__5517\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22408\
        );

    \I__5516\ : CascadeMux
    port map (
            O => \N__22420\,
            I => \N__22403\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__22417\,
            I => \N__22399\
        );

    \I__5514\ : InMux
    port map (
            O => \N__22416\,
            I => \N__22396\
        );

    \I__5513\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22393\
        );

    \I__5512\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22390\
        );

    \I__5511\ : InMux
    port map (
            O => \N__22411\,
            I => \N__22387\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__22408\,
            I => \N__22384\
        );

    \I__5509\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22379\
        );

    \I__5508\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22379\
        );

    \I__5507\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22373\
        );

    \I__5506\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22373\
        );

    \I__5505\ : Span12Mux_s3_h
    port map (
            O => \N__22399\,
            I => \N__22370\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__22396\,
            I => \N__22365\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22365\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__22390\,
            I => \N__22360\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__22387\,
            I => \N__22360\
        );

    \I__5500\ : Span4Mux_s3_h
    port map (
            O => \N__22384\,
            I => \N__22355\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__22379\,
            I => \N__22355\
        );

    \I__5498\ : InMux
    port map (
            O => \N__22378\,
            I => \N__22352\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__22373\,
            I => \Lab_UT.state_i_3_2_rep2\
        );

    \I__5496\ : Odrv12
    port map (
            O => \N__22370\,
            I => \Lab_UT.state_i_3_2_rep2\
        );

    \I__5495\ : Odrv12
    port map (
            O => \N__22365\,
            I => \Lab_UT.state_i_3_2_rep2\
        );

    \I__5494\ : Odrv4
    port map (
            O => \N__22360\,
            I => \Lab_UT.state_i_3_2_rep2\
        );

    \I__5493\ : Odrv4
    port map (
            O => \N__22355\,
            I => \Lab_UT.state_i_3_2_rep2\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__22352\,
            I => \Lab_UT.state_i_3_2_rep2\
        );

    \I__5491\ : CascadeMux
    port map (
            O => \N__22339\,
            I => \N__22336\
        );

    \I__5490\ : InMux
    port map (
            O => \N__22336\,
            I => \N__22328\
        );

    \I__5489\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22320\
        );

    \I__5488\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22316\
        );

    \I__5487\ : CascadeMux
    port map (
            O => \N__22333\,
            I => \N__22313\
        );

    \I__5486\ : CascadeMux
    port map (
            O => \N__22332\,
            I => \N__22309\
        );

    \I__5485\ : CascadeMux
    port map (
            O => \N__22331\,
            I => \N__22306\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__22328\,
            I => \N__22298\
        );

    \I__5483\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22293\
        );

    \I__5482\ : InMux
    port map (
            O => \N__22326\,
            I => \N__22284\
        );

    \I__5481\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22284\
        );

    \I__5480\ : InMux
    port map (
            O => \N__22324\,
            I => \N__22284\
        );

    \I__5479\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22284\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__22320\,
            I => \N__22281\
        );

    \I__5477\ : InMux
    port map (
            O => \N__22319\,
            I => \N__22278\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__22316\,
            I => \N__22275\
        );

    \I__5475\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22270\
        );

    \I__5474\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22270\
        );

    \I__5473\ : InMux
    port map (
            O => \N__22309\,
            I => \N__22263\
        );

    \I__5472\ : InMux
    port map (
            O => \N__22306\,
            I => \N__22263\
        );

    \I__5471\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22260\
        );

    \I__5470\ : CascadeMux
    port map (
            O => \N__22304\,
            I => \N__22254\
        );

    \I__5469\ : InMux
    port map (
            O => \N__22303\,
            I => \N__22248\
        );

    \I__5468\ : InMux
    port map (
            O => \N__22302\,
            I => \N__22248\
        );

    \I__5467\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22245\
        );

    \I__5466\ : Span4Mux_v
    port map (
            O => \N__22298\,
            I => \N__22242\
        );

    \I__5465\ : InMux
    port map (
            O => \N__22297\,
            I => \N__22239\
        );

    \I__5464\ : InMux
    port map (
            O => \N__22296\,
            I => \N__22236\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__22293\,
            I => \N__22231\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__22284\,
            I => \N__22231\
        );

    \I__5461\ : Span4Mux_s3_v
    port map (
            O => \N__22281\,
            I => \N__22226\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__22278\,
            I => \N__22226\
        );

    \I__5459\ : Span4Mux_s3_v
    port map (
            O => \N__22275\,
            I => \N__22221\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22221\
        );

    \I__5457\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22216\
        );

    \I__5456\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22216\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__22263\,
            I => \N__22213\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__22260\,
            I => \N__22210\
        );

    \I__5453\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22207\
        );

    \I__5452\ : InMux
    port map (
            O => \N__22258\,
            I => \N__22202\
        );

    \I__5451\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22202\
        );

    \I__5450\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22199\
        );

    \I__5449\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22196\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__22248\,
            I => \N__22193\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__22245\,
            I => \N__22187\
        );

    \I__5446\ : Span4Mux_v
    port map (
            O => \N__22242\,
            I => \N__22184\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__22239\,
            I => \N__22177\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__22236\,
            I => \N__22177\
        );

    \I__5443\ : Span4Mux_v
    port map (
            O => \N__22231\,
            I => \N__22177\
        );

    \I__5442\ : Span4Mux_v
    port map (
            O => \N__22226\,
            I => \N__22172\
        );

    \I__5441\ : Span4Mux_v
    port map (
            O => \N__22221\,
            I => \N__22172\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__22216\,
            I => \N__22169\
        );

    \I__5439\ : Span4Mux_s2_h
    port map (
            O => \N__22213\,
            I => \N__22160\
        );

    \I__5438\ : Span4Mux_h
    port map (
            O => \N__22210\,
            I => \N__22160\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__22207\,
            I => \N__22160\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__22202\,
            I => \N__22160\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__22199\,
            I => \N__22153\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__22196\,
            I => \N__22153\
        );

    \I__5433\ : Span4Mux_v
    port map (
            O => \N__22193\,
            I => \N__22153\
        );

    \I__5432\ : CascadeMux
    port map (
            O => \N__22192\,
            I => \N__22149\
        );

    \I__5431\ : CascadeMux
    port map (
            O => \N__22191\,
            I => \N__22146\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__22190\,
            I => \N__22143\
        );

    \I__5429\ : Span4Mux_s2_h
    port map (
            O => \N__22187\,
            I => \N__22140\
        );

    \I__5428\ : Span4Mux_v
    port map (
            O => \N__22184\,
            I => \N__22135\
        );

    \I__5427\ : Span4Mux_v
    port map (
            O => \N__22177\,
            I => \N__22135\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__22172\,
            I => \N__22130\
        );

    \I__5425\ : Span4Mux_h
    port map (
            O => \N__22169\,
            I => \N__22130\
        );

    \I__5424\ : Span4Mux_v
    port map (
            O => \N__22160\,
            I => \N__22125\
        );

    \I__5423\ : Span4Mux_h
    port map (
            O => \N__22153\,
            I => \N__22125\
        );

    \I__5422\ : InMux
    port map (
            O => \N__22152\,
            I => \N__22120\
        );

    \I__5421\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22120\
        );

    \I__5420\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22115\
        );

    \I__5419\ : InMux
    port map (
            O => \N__22143\,
            I => \N__22115\
        );

    \I__5418\ : Odrv4
    port map (
            O => \N__22140\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__5417\ : Odrv4
    port map (
            O => \N__22135\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__5416\ : Odrv4
    port map (
            O => \N__22130\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__5415\ : Odrv4
    port map (
            O => \N__22125\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__22120\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__22115\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__5412\ : CascadeMux
    port map (
            O => \N__22102\,
            I => \N__22097\
        );

    \I__5411\ : CascadeMux
    port map (
            O => \N__22101\,
            I => \N__22087\
        );

    \I__5410\ : CascadeMux
    port map (
            O => \N__22100\,
            I => \N__22084\
        );

    \I__5409\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22081\
        );

    \I__5408\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22078\
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__22095\,
            I => \N__22074\
        );

    \I__5406\ : CascadeMux
    port map (
            O => \N__22094\,
            I => \N__22070\
        );

    \I__5405\ : CascadeMux
    port map (
            O => \N__22093\,
            I => \N__22066\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__22092\,
            I => \N__22062\
        );

    \I__5403\ : CascadeMux
    port map (
            O => \N__22091\,
            I => \N__22059\
        );

    \I__5402\ : InMux
    port map (
            O => \N__22090\,
            I => \N__22056\
        );

    \I__5401\ : InMux
    port map (
            O => \N__22087\,
            I => \N__22051\
        );

    \I__5400\ : InMux
    port map (
            O => \N__22084\,
            I => \N__22051\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__22081\,
            I => \N__22046\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__22078\,
            I => \N__22046\
        );

    \I__5397\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22041\
        );

    \I__5396\ : InMux
    port map (
            O => \N__22074\,
            I => \N__22041\
        );

    \I__5395\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22036\
        );

    \I__5394\ : InMux
    port map (
            O => \N__22070\,
            I => \N__22036\
        );

    \I__5393\ : CascadeMux
    port map (
            O => \N__22069\,
            I => \N__22033\
        );

    \I__5392\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22030\
        );

    \I__5391\ : CascadeMux
    port map (
            O => \N__22065\,
            I => \N__22027\
        );

    \I__5390\ : InMux
    port map (
            O => \N__22062\,
            I => \N__22024\
        );

    \I__5389\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22021\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__22056\,
            I => \N__22014\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__22051\,
            I => \N__22014\
        );

    \I__5386\ : Span4Mux_v
    port map (
            O => \N__22046\,
            I => \N__22014\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__22041\,
            I => \N__22009\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__22036\,
            I => \N__22009\
        );

    \I__5383\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22006\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__22030\,
            I => \N__22003\
        );

    \I__5381\ : InMux
    port map (
            O => \N__22027\,
            I => \N__22000\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__22024\,
            I => \N__21997\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__22021\,
            I => \N__21990\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__22014\,
            I => \N__21990\
        );

    \I__5377\ : Span4Mux_v
    port map (
            O => \N__22009\,
            I => \N__21990\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__22006\,
            I => \N__21985\
        );

    \I__5375\ : Span4Mux_h
    port map (
            O => \N__22003\,
            I => \N__21985\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__22000\,
            I => \Lab_UT.scctrl.state_i_3_0_rep2\
        );

    \I__5373\ : Odrv12
    port map (
            O => \N__21997\,
            I => \Lab_UT.scctrl.state_i_3_0_rep2\
        );

    \I__5372\ : Odrv4
    port map (
            O => \N__21990\,
            I => \Lab_UT.scctrl.state_i_3_0_rep2\
        );

    \I__5371\ : Odrv4
    port map (
            O => \N__21985\,
            I => \Lab_UT.scctrl.state_i_3_0_rep2\
        );

    \I__5370\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21972\
        );

    \I__5369\ : InMux
    port map (
            O => \N__21975\,
            I => \N__21969\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__21972\,
            I => \N__21964\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__21969\,
            I => \N__21964\
        );

    \I__5366\ : Odrv4
    port map (
            O => \N__21964\,
            I => rst_i_3_fast
        );

    \I__5365\ : InMux
    port map (
            O => \N__21961\,
            I => \N__21958\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__21958\,
            I => \Lab_UT.scctrl.g1_i_0\
        );

    \I__5363\ : InMux
    port map (
            O => \N__21955\,
            I => \N__21952\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__21952\,
            I => \N__21944\
        );

    \I__5361\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21938\
        );

    \I__5360\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21933\
        );

    \I__5359\ : InMux
    port map (
            O => \N__21949\,
            I => \N__21933\
        );

    \I__5358\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21930\
        );

    \I__5357\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21924\
        );

    \I__5356\ : Span4Mux_s1_v
    port map (
            O => \N__21944\,
            I => \N__21919\
        );

    \I__5355\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21916\
        );

    \I__5354\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21913\
        );

    \I__5353\ : InMux
    port map (
            O => \N__21941\,
            I => \N__21910\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__21938\,
            I => \N__21907\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__21933\,
            I => \N__21904\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__21930\,
            I => \N__21901\
        );

    \I__5349\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21896\
        );

    \I__5348\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21896\
        );

    \I__5347\ : InMux
    port map (
            O => \N__21927\,
            I => \N__21893\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__21924\,
            I => \N__21890\
        );

    \I__5345\ : InMux
    port map (
            O => \N__21923\,
            I => \N__21887\
        );

    \I__5344\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21884\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__21919\,
            I => \N__21879\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__21916\,
            I => \N__21879\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__21913\,
            I => \N__21874\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__21910\,
            I => \N__21874\
        );

    \I__5339\ : Span4Mux_v
    port map (
            O => \N__21907\,
            I => \N__21871\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__21904\,
            I => \N__21862\
        );

    \I__5337\ : Span4Mux_s2_h
    port map (
            O => \N__21901\,
            I => \N__21862\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__21896\,
            I => \N__21859\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__21893\,
            I => \N__21856\
        );

    \I__5334\ : Span12Mux_s11_h
    port map (
            O => \N__21890\,
            I => \N__21853\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__21887\,
            I => \N__21850\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__21884\,
            I => \N__21843\
        );

    \I__5331\ : Span4Mux_v
    port map (
            O => \N__21879\,
            I => \N__21843\
        );

    \I__5330\ : Span4Mux_h
    port map (
            O => \N__21874\,
            I => \N__21843\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__21871\,
            I => \N__21840\
        );

    \I__5328\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21837\
        );

    \I__5327\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21830\
        );

    \I__5326\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21830\
        );

    \I__5325\ : InMux
    port map (
            O => \N__21867\,
            I => \N__21830\
        );

    \I__5324\ : Span4Mux_v
    port map (
            O => \N__21862\,
            I => \N__21823\
        );

    \I__5323\ : Span4Mux_s2_h
    port map (
            O => \N__21859\,
            I => \N__21823\
        );

    \I__5322\ : Span4Mux_h
    port map (
            O => \N__21856\,
            I => \N__21823\
        );

    \I__5321\ : Span12Mux_v
    port map (
            O => \N__21853\,
            I => \N__21820\
        );

    \I__5320\ : Span4Mux_s2_h
    port map (
            O => \N__21850\,
            I => \N__21815\
        );

    \I__5319\ : Span4Mux_v
    port map (
            O => \N__21843\,
            I => \N__21815\
        );

    \I__5318\ : Odrv4
    port map (
            O => \N__21840\,
            I => \Lab_UT.state_i_3_0\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__21837\,
            I => \Lab_UT.state_i_3_0\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__21830\,
            I => \Lab_UT.state_i_3_0\
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__21823\,
            I => \Lab_UT.state_i_3_0\
        );

    \I__5314\ : Odrv12
    port map (
            O => \N__21820\,
            I => \Lab_UT.state_i_3_0\
        );

    \I__5313\ : Odrv4
    port map (
            O => \N__21815\,
            I => \Lab_UT.state_i_3_0\
        );

    \I__5312\ : CascadeMux
    port map (
            O => \N__21802\,
            I => \N__21799\
        );

    \I__5311\ : InMux
    port map (
            O => \N__21799\,
            I => \N__21796\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__21796\,
            I => \Lab_UT.scctrl.g0_0_i_a8_3_1\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__21793\,
            I => \N__21784\
        );

    \I__5308\ : CascadeMux
    port map (
            O => \N__21792\,
            I => \N__21779\
        );

    \I__5307\ : CascadeMux
    port map (
            O => \N__21791\,
            I => \N__21776\
        );

    \I__5306\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21771\
        );

    \I__5305\ : InMux
    port map (
            O => \N__21789\,
            I => \N__21771\
        );

    \I__5304\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21757\
        );

    \I__5303\ : InMux
    port map (
            O => \N__21787\,
            I => \N__21753\
        );

    \I__5302\ : InMux
    port map (
            O => \N__21784\,
            I => \N__21750\
        );

    \I__5301\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21747\
        );

    \I__5300\ : CascadeMux
    port map (
            O => \N__21782\,
            I => \N__21744\
        );

    \I__5299\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21739\
        );

    \I__5298\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21736\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__21771\,
            I => \N__21732\
        );

    \I__5296\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21729\
        );

    \I__5295\ : InMux
    port map (
            O => \N__21769\,
            I => \N__21726\
        );

    \I__5294\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21723\
        );

    \I__5293\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21716\
        );

    \I__5292\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21716\
        );

    \I__5291\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21716\
        );

    \I__5290\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21707\
        );

    \I__5289\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21707\
        );

    \I__5288\ : InMux
    port map (
            O => \N__21762\,
            I => \N__21707\
        );

    \I__5287\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21702\
        );

    \I__5286\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21702\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__21757\,
            I => \N__21699\
        );

    \I__5284\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21695\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__21753\,
            I => \N__21692\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__21750\,
            I => \N__21689\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__21747\,
            I => \N__21685\
        );

    \I__5280\ : InMux
    port map (
            O => \N__21744\,
            I => \N__21682\
        );

    \I__5279\ : InMux
    port map (
            O => \N__21743\,
            I => \N__21677\
        );

    \I__5278\ : InMux
    port map (
            O => \N__21742\,
            I => \N__21677\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__21739\,
            I => \N__21674\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__21736\,
            I => \N__21670\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__21735\,
            I => \N__21665\
        );

    \I__5274\ : Span4Mux_v
    port map (
            O => \N__21732\,
            I => \N__21662\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__21729\,
            I => \N__21659\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__21726\,
            I => \N__21656\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__21723\,
            I => \N__21651\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21651\
        );

    \I__5269\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21646\
        );

    \I__5268\ : InMux
    port map (
            O => \N__21714\,
            I => \N__21646\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__21707\,
            I => \N__21641\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__21702\,
            I => \N__21641\
        );

    \I__5265\ : Span4Mux_h
    port map (
            O => \N__21699\,
            I => \N__21638\
        );

    \I__5264\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21635\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__21695\,
            I => \N__21628\
        );

    \I__5262\ : Span4Mux_v
    port map (
            O => \N__21692\,
            I => \N__21628\
        );

    \I__5261\ : Span4Mux_s1_h
    port map (
            O => \N__21689\,
            I => \N__21628\
        );

    \I__5260\ : InMux
    port map (
            O => \N__21688\,
            I => \N__21625\
        );

    \I__5259\ : Span12Mux_s5_h
    port map (
            O => \N__21685\,
            I => \N__21618\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__21682\,
            I => \N__21618\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__21677\,
            I => \N__21618\
        );

    \I__5256\ : Span4Mux_v
    port map (
            O => \N__21674\,
            I => \N__21615\
        );

    \I__5255\ : InMux
    port map (
            O => \N__21673\,
            I => \N__21612\
        );

    \I__5254\ : Span4Mux_v
    port map (
            O => \N__21670\,
            I => \N__21609\
        );

    \I__5253\ : InMux
    port map (
            O => \N__21669\,
            I => \N__21602\
        );

    \I__5252\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21602\
        );

    \I__5251\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21602\
        );

    \I__5250\ : Span4Mux_h
    port map (
            O => \N__21662\,
            I => \N__21593\
        );

    \I__5249\ : Span4Mux_h
    port map (
            O => \N__21659\,
            I => \N__21593\
        );

    \I__5248\ : Span4Mux_h
    port map (
            O => \N__21656\,
            I => \N__21593\
        );

    \I__5247\ : Span4Mux_v
    port map (
            O => \N__21651\,
            I => \N__21593\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__21646\,
            I => \N__21588\
        );

    \I__5245\ : Span4Mux_v
    port map (
            O => \N__21641\,
            I => \N__21588\
        );

    \I__5244\ : Span4Mux_v
    port map (
            O => \N__21638\,
            I => \N__21581\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__21635\,
            I => \N__21581\
        );

    \I__5242\ : Span4Mux_h
    port map (
            O => \N__21628\,
            I => \N__21581\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__21625\,
            I => \Lab_UT.state_1\
        );

    \I__5240\ : Odrv12
    port map (
            O => \N__21618\,
            I => \Lab_UT.state_1\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__21615\,
            I => \Lab_UT.state_1\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__21612\,
            I => \Lab_UT.state_1\
        );

    \I__5237\ : Odrv4
    port map (
            O => \N__21609\,
            I => \Lab_UT.state_1\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__21602\,
            I => \Lab_UT.state_1\
        );

    \I__5235\ : Odrv4
    port map (
            O => \N__21593\,
            I => \Lab_UT.state_1\
        );

    \I__5234\ : Odrv4
    port map (
            O => \N__21588\,
            I => \Lab_UT.state_1\
        );

    \I__5233\ : Odrv4
    port map (
            O => \N__21581\,
            I => \Lab_UT.state_1\
        );

    \I__5232\ : InMux
    port map (
            O => \N__21562\,
            I => \N__21559\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__21559\,
            I => \Lab_UT.scctrl.state_1_RNO_3Z0Z_0\
        );

    \I__5230\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21553\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__21553\,
            I => \N__21550\
        );

    \I__5228\ : Odrv4
    port map (
            O => \N__21550\,
            I => \Lab_UT.scctrl.N_13_0\
        );

    \I__5227\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21543\
        );

    \I__5226\ : InMux
    port map (
            O => \N__21546\,
            I => \N__21540\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__21543\,
            I => \N__21537\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__21540\,
            I => \N__21534\
        );

    \I__5223\ : Span4Mux_s0_h
    port map (
            O => \N__21537\,
            I => \N__21531\
        );

    \I__5222\ : Span4Mux_h
    port map (
            O => \N__21534\,
            I => \N__21525\
        );

    \I__5221\ : Span4Mux_h
    port map (
            O => \N__21531\,
            I => \N__21522\
        );

    \I__5220\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21515\
        );

    \I__5219\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21515\
        );

    \I__5218\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21515\
        );

    \I__5217\ : Odrv4
    port map (
            O => \N__21525\,
            I => \Lab_UT.N_191\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__21522\,
            I => \Lab_UT.N_191\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__21515\,
            I => \Lab_UT.N_191\
        );

    \I__5214\ : CascadeMux
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__5213\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21502\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__21502\,
            I => \N__21499\
        );

    \I__5211\ : Span4Mux_s1_h
    port map (
            O => \N__21499\,
            I => \N__21496\
        );

    \I__5210\ : Span4Mux_h
    port map (
            O => \N__21496\,
            I => \N__21493\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__21493\,
            I => \Lab_UT.scctrl.G_24_i_a4_0_1\
        );

    \I__5208\ : InMux
    port map (
            O => \N__21490\,
            I => \N__21486\
        );

    \I__5207\ : InMux
    port map (
            O => \N__21489\,
            I => \N__21483\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__21486\,
            I => \N__21480\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__21483\,
            I => \N__21474\
        );

    \I__5204\ : Span4Mux_v
    port map (
            O => \N__21480\,
            I => \N__21471\
        );

    \I__5203\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21464\
        );

    \I__5202\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21464\
        );

    \I__5201\ : InMux
    port map (
            O => \N__21477\,
            I => \N__21464\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__21474\,
            I => \N__21457\
        );

    \I__5199\ : Span4Mux_h
    port map (
            O => \N__21471\,
            I => \N__21457\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__21464\,
            I => \N__21457\
        );

    \I__5197\ : Odrv4
    port map (
            O => \N__21457\,
            I => \Lab_UT.next_state_1_0_0_3\
        );

    \I__5196\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21451\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__21451\,
            I => \N__21448\
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__21448\,
            I => \Lab_UT.scctrl.N_10_2\
        );

    \I__5193\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21441\
        );

    \I__5192\ : CascadeMux
    port map (
            O => \N__21444\,
            I => \N__21436\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__21441\,
            I => \N__21433\
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__21440\,
            I => \N__21429\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__21439\,
            I => \N__21421\
        );

    \I__5188\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21416\
        );

    \I__5187\ : Span4Mux_v
    port map (
            O => \N__21433\,
            I => \N__21413\
        );

    \I__5186\ : InMux
    port map (
            O => \N__21432\,
            I => \N__21410\
        );

    \I__5185\ : InMux
    port map (
            O => \N__21429\,
            I => \N__21402\
        );

    \I__5184\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21402\
        );

    \I__5183\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21392\
        );

    \I__5182\ : InMux
    port map (
            O => \N__21426\,
            I => \N__21392\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__21425\,
            I => \N__21389\
        );

    \I__5180\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21383\
        );

    \I__5179\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21383\
        );

    \I__5178\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21378\
        );

    \I__5177\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21378\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__21416\,
            I => \N__21369\
        );

    \I__5175\ : Span4Mux_v
    port map (
            O => \N__21413\,
            I => \N__21369\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__21410\,
            I => \N__21369\
        );

    \I__5173\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21364\
        );

    \I__5172\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21364\
        );

    \I__5171\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21359\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__21402\,
            I => \N__21356\
        );

    \I__5169\ : InMux
    port map (
            O => \N__21401\,
            I => \N__21351\
        );

    \I__5168\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21351\
        );

    \I__5167\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21344\
        );

    \I__5166\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21344\
        );

    \I__5165\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21344\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21341\
        );

    \I__5163\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21336\
        );

    \I__5162\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21336\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__21383\,
            I => \N__21331\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__21378\,
            I => \N__21331\
        );

    \I__5159\ : InMux
    port map (
            O => \N__21377\,
            I => \N__21328\
        );

    \I__5158\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21325\
        );

    \I__5157\ : Span4Mux_v
    port map (
            O => \N__21369\,
            I => \N__21321\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__21364\,
            I => \N__21318\
        );

    \I__5155\ : InMux
    port map (
            O => \N__21363\,
            I => \N__21313\
        );

    \I__5154\ : InMux
    port map (
            O => \N__21362\,
            I => \N__21313\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__21359\,
            I => \N__21306\
        );

    \I__5152\ : Span4Mux_h
    port map (
            O => \N__21356\,
            I => \N__21306\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__21351\,
            I => \N__21306\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__21344\,
            I => \N__21303\
        );

    \I__5149\ : Span4Mux_v
    port map (
            O => \N__21341\,
            I => \N__21300\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__21336\,
            I => \N__21291\
        );

    \I__5147\ : Span4Mux_v
    port map (
            O => \N__21331\,
            I => \N__21291\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__21328\,
            I => \N__21291\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__21325\,
            I => \N__21291\
        );

    \I__5144\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21287\
        );

    \I__5143\ : Span4Mux_v
    port map (
            O => \N__21321\,
            I => \N__21284\
        );

    \I__5142\ : Span4Mux_h
    port map (
            O => \N__21318\,
            I => \N__21277\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__21313\,
            I => \N__21277\
        );

    \I__5140\ : Span4Mux_h
    port map (
            O => \N__21306\,
            I => \N__21277\
        );

    \I__5139\ : Span4Mux_h
    port map (
            O => \N__21303\,
            I => \N__21272\
        );

    \I__5138\ : Span4Mux_h
    port map (
            O => \N__21300\,
            I => \N__21272\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__21291\,
            I => \N__21269\
        );

    \I__5136\ : InMux
    port map (
            O => \N__21290\,
            I => \N__21266\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__21287\,
            I => \Lab_UT.N_169_0\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__21284\,
            I => \Lab_UT.N_169_0\
        );

    \I__5133\ : Odrv4
    port map (
            O => \N__21277\,
            I => \Lab_UT.N_169_0\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__21272\,
            I => \Lab_UT.N_169_0\
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__21269\,
            I => \Lab_UT.N_169_0\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__21266\,
            I => \Lab_UT.N_169_0\
        );

    \I__5129\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21250\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__21250\,
            I => \N__21245\
        );

    \I__5127\ : InMux
    port map (
            O => \N__21249\,
            I => \N__21242\
        );

    \I__5126\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21239\
        );

    \I__5125\ : Span4Mux_v
    port map (
            O => \N__21245\,
            I => \N__21236\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__21242\,
            I => \N__21233\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__21239\,
            I => \N__21230\
        );

    \I__5122\ : Span4Mux_v
    port map (
            O => \N__21236\,
            I => \N__21227\
        );

    \I__5121\ : Span12Mux_v
    port map (
            O => \N__21233\,
            I => \N__21224\
        );

    \I__5120\ : Span4Mux_h
    port map (
            O => \N__21230\,
            I => \N__21221\
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__21227\,
            I => \Lab_UT.scctrl.N_223_1\
        );

    \I__5118\ : Odrv12
    port map (
            O => \N__21224\,
            I => \Lab_UT.scctrl.N_223_1\
        );

    \I__5117\ : Odrv4
    port map (
            O => \N__21221\,
            I => \Lab_UT.scctrl.N_223_1\
        );

    \I__5116\ : IoInMux
    port map (
            O => \N__21214\,
            I => \N__21211\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__21211\,
            I => led_c_4
        );

    \I__5114\ : CascadeMux
    port map (
            O => \N__21208\,
            I => \N__21203\
        );

    \I__5113\ : CascadeMux
    port map (
            O => \N__21207\,
            I => \N__21197\
        );

    \I__5112\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21192\
        );

    \I__5111\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21186\
        );

    \I__5110\ : CascadeMux
    port map (
            O => \N__21202\,
            I => \N__21182\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__21201\,
            I => \N__21179\
        );

    \I__5108\ : CascadeMux
    port map (
            O => \N__21200\,
            I => \N__21176\
        );

    \I__5107\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21169\
        );

    \I__5106\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21166\
        );

    \I__5105\ : CascadeMux
    port map (
            O => \N__21195\,
            I => \N__21162\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__21192\,
            I => \N__21157\
        );

    \I__5103\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21152\
        );

    \I__5102\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21152\
        );

    \I__5101\ : InMux
    port map (
            O => \N__21189\,
            I => \N__21149\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21186\,
            I => \N__21146\
        );

    \I__5099\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21143\
        );

    \I__5098\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21138\
        );

    \I__5097\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21138\
        );

    \I__5096\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21135\
        );

    \I__5095\ : InMux
    port map (
            O => \N__21175\,
            I => \N__21130\
        );

    \I__5094\ : InMux
    port map (
            O => \N__21174\,
            I => \N__21130\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__21173\,
            I => \N__21123\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__21172\,
            I => \N__21120\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__21169\,
            I => \N__21117\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__21166\,
            I => \N__21114\
        );

    \I__5089\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21109\
        );

    \I__5088\ : InMux
    port map (
            O => \N__21162\,
            I => \N__21109\
        );

    \I__5087\ : InMux
    port map (
            O => \N__21161\,
            I => \N__21104\
        );

    \I__5086\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21104\
        );

    \I__5085\ : Span4Mux_s3_h
    port map (
            O => \N__21157\,
            I => \N__21095\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__21152\,
            I => \N__21095\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__21149\,
            I => \N__21095\
        );

    \I__5082\ : Span4Mux_h
    port map (
            O => \N__21146\,
            I => \N__21095\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__21143\,
            I => \N__21092\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__21138\,
            I => \N__21087\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__21135\,
            I => \N__21087\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__21130\,
            I => \N__21084\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__21129\,
            I => \N__21081\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__21128\,
            I => \N__21078\
        );

    \I__5075\ : InMux
    port map (
            O => \N__21127\,
            I => \N__21075\
        );

    \I__5074\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21072\
        );

    \I__5073\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21069\
        );

    \I__5072\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21066\
        );

    \I__5071\ : Span12Mux_s4_h
    port map (
            O => \N__21117\,
            I => \N__21059\
        );

    \I__5070\ : Span12Mux_s8_v
    port map (
            O => \N__21114\,
            I => \N__21059\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__21109\,
            I => \N__21059\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__21104\,
            I => \N__21054\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__21095\,
            I => \N__21054\
        );

    \I__5066\ : Span4Mux_v
    port map (
            O => \N__21092\,
            I => \N__21047\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__21087\,
            I => \N__21047\
        );

    \I__5064\ : Span4Mux_v
    port map (
            O => \N__21084\,
            I => \N__21047\
        );

    \I__5063\ : InMux
    port map (
            O => \N__21081\,
            I => \N__21042\
        );

    \I__5062\ : InMux
    port map (
            O => \N__21078\,
            I => \N__21042\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__21075\,
            I => \Lab_UT.un1_state_3_1\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__21072\,
            I => \Lab_UT.un1_state_3_1\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__21069\,
            I => \Lab_UT.un1_state_3_1\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__21066\,
            I => \Lab_UT.un1_state_3_1\
        );

    \I__5057\ : Odrv12
    port map (
            O => \N__21059\,
            I => \Lab_UT.un1_state_3_1\
        );

    \I__5056\ : Odrv4
    port map (
            O => \N__21054\,
            I => \Lab_UT.un1_state_3_1\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__21047\,
            I => \Lab_UT.un1_state_3_1\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__21042\,
            I => \Lab_UT.un1_state_3_1\
        );

    \I__5053\ : InMux
    port map (
            O => \N__21025\,
            I => \N__21016\
        );

    \I__5052\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21008\
        );

    \I__5051\ : InMux
    port map (
            O => \N__21023\,
            I => \N__21003\
        );

    \I__5050\ : InMux
    port map (
            O => \N__21022\,
            I => \N__21000\
        );

    \I__5049\ : InMux
    port map (
            O => \N__21021\,
            I => \N__20997\
        );

    \I__5048\ : InMux
    port map (
            O => \N__21020\,
            I => \N__20992\
        );

    \I__5047\ : InMux
    port map (
            O => \N__21019\,
            I => \N__20992\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__21016\,
            I => \N__20978\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21015\,
            I => \N__20975\
        );

    \I__5044\ : InMux
    port map (
            O => \N__21014\,
            I => \N__20972\
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__21013\,
            I => \N__20969\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21012\,
            I => \N__20964\
        );

    \I__5041\ : InMux
    port map (
            O => \N__21011\,
            I => \N__20964\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__21008\,
            I => \N__20961\
        );

    \I__5039\ : InMux
    port map (
            O => \N__21007\,
            I => \N__20956\
        );

    \I__5038\ : InMux
    port map (
            O => \N__21006\,
            I => \N__20956\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__21003\,
            I => \N__20953\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__21000\,
            I => \N__20948\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__20997\,
            I => \N__20948\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__20992\,
            I => \N__20945\
        );

    \I__5033\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20940\
        );

    \I__5032\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20940\
        );

    \I__5031\ : InMux
    port map (
            O => \N__20989\,
            I => \N__20937\
        );

    \I__5030\ : InMux
    port map (
            O => \N__20988\,
            I => \N__20932\
        );

    \I__5029\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20932\
        );

    \I__5028\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20920\
        );

    \I__5027\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20920\
        );

    \I__5026\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20920\
        );

    \I__5025\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20913\
        );

    \I__5024\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20913\
        );

    \I__5023\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20913\
        );

    \I__5022\ : Span4Mux_s1_h
    port map (
            O => \N__20978\,
            I => \N__20905\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20905\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__20972\,
            I => \N__20902\
        );

    \I__5019\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20899\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__20964\,
            I => \N__20892\
        );

    \I__5017\ : Span4Mux_h
    port map (
            O => \N__20961\,
            I => \N__20892\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__20956\,
            I => \N__20892\
        );

    \I__5015\ : Span4Mux_v
    port map (
            O => \N__20953\,
            I => \N__20883\
        );

    \I__5014\ : Span4Mux_v
    port map (
            O => \N__20948\,
            I => \N__20883\
        );

    \I__5013\ : Span4Mux_h
    port map (
            O => \N__20945\,
            I => \N__20883\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__20940\,
            I => \N__20883\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__20937\,
            I => \N__20878\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__20932\,
            I => \N__20878\
        );

    \I__5009\ : InMux
    port map (
            O => \N__20931\,
            I => \N__20871\
        );

    \I__5008\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20871\
        );

    \I__5007\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20871\
        );

    \I__5006\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20866\
        );

    \I__5005\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20866\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__20920\,
            I => \N__20861\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__20913\,
            I => \N__20861\
        );

    \I__5002\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20854\
        );

    \I__5001\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20854\
        );

    \I__5000\ : InMux
    port map (
            O => \N__20910\,
            I => \N__20854\
        );

    \I__4999\ : Span4Mux_h
    port map (
            O => \N__20905\,
            I => \N__20847\
        );

    \I__4998\ : Span4Mux_v
    port map (
            O => \N__20902\,
            I => \N__20847\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__20899\,
            I => \N__20847\
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__20892\,
            I => \L4_PrintBuf\
        );

    \I__4995\ : Odrv4
    port map (
            O => \N__20883\,
            I => \L4_PrintBuf\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__20878\,
            I => \L4_PrintBuf\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__20871\,
            I => \L4_PrintBuf\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__20866\,
            I => \L4_PrintBuf\
        );

    \I__4991\ : Odrv12
    port map (
            O => \N__20861\,
            I => \L4_PrintBuf\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__20854\,
            I => \L4_PrintBuf\
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__20847\,
            I => \L4_PrintBuf\
        );

    \I__4988\ : InMux
    port map (
            O => \N__20830\,
            I => \N__20827\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__20827\,
            I => \N__20824\
        );

    \I__4986\ : Span4Mux_h
    port map (
            O => \N__20824\,
            I => \N__20821\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__20821\,
            I => \Lab_UT.scctrl.m26_i_o4_1_2\
        );

    \I__4984\ : CascadeMux
    port map (
            O => \N__20818\,
            I => \Lab_UT.scctrl.G_24_i_o3_0_0_cascade_\
        );

    \I__4983\ : CascadeMux
    port map (
            O => \N__20815\,
            I => \N__20811\
        );

    \I__4982\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20800\
        );

    \I__4981\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20797\
        );

    \I__4980\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20792\
        );

    \I__4979\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20792\
        );

    \I__4978\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20788\
        );

    \I__4977\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20781\
        );

    \I__4976\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20776\
        );

    \I__4975\ : InMux
    port map (
            O => \N__20805\,
            I => \N__20776\
        );

    \I__4974\ : InMux
    port map (
            O => \N__20804\,
            I => \N__20771\
        );

    \I__4973\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20771\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__20800\,
            I => \N__20768\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__20797\,
            I => \N__20765\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__20792\,
            I => \N__20762\
        );

    \I__4969\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20759\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__20788\,
            I => \N__20754\
        );

    \I__4967\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20749\
        );

    \I__4966\ : InMux
    port map (
            O => \N__20786\,
            I => \N__20742\
        );

    \I__4965\ : InMux
    port map (
            O => \N__20785\,
            I => \N__20742\
        );

    \I__4964\ : InMux
    port map (
            O => \N__20784\,
            I => \N__20742\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__20781\,
            I => \N__20737\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__20776\,
            I => \N__20737\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__20771\,
            I => \N__20734\
        );

    \I__4960\ : Span4Mux_s1_h
    port map (
            O => \N__20768\,
            I => \N__20729\
        );

    \I__4959\ : Span4Mux_v
    port map (
            O => \N__20765\,
            I => \N__20729\
        );

    \I__4958\ : Span4Mux_v
    port map (
            O => \N__20762\,
            I => \N__20726\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__20759\,
            I => \N__20723\
        );

    \I__4956\ : InMux
    port map (
            O => \N__20758\,
            I => \N__20720\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__20757\,
            I => \N__20714\
        );

    \I__4954\ : Span4Mux_v
    port map (
            O => \N__20754\,
            I => \N__20710\
        );

    \I__4953\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20707\
        );

    \I__4952\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20704\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__20749\,
            I => \N__20697\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__20742\,
            I => \N__20697\
        );

    \I__4949\ : Span4Mux_h
    port map (
            O => \N__20737\,
            I => \N__20697\
        );

    \I__4948\ : Span4Mux_v
    port map (
            O => \N__20734\,
            I => \N__20692\
        );

    \I__4947\ : Span4Mux_h
    port map (
            O => \N__20729\,
            I => \N__20692\
        );

    \I__4946\ : Span4Mux_h
    port map (
            O => \N__20726\,
            I => \N__20685\
        );

    \I__4945\ : Span4Mux_v
    port map (
            O => \N__20723\,
            I => \N__20685\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__20720\,
            I => \N__20685\
        );

    \I__4943\ : InMux
    port map (
            O => \N__20719\,
            I => \N__20682\
        );

    \I__4942\ : InMux
    port map (
            O => \N__20718\,
            I => \N__20679\
        );

    \I__4941\ : InMux
    port map (
            O => \N__20717\,
            I => \N__20676\
        );

    \I__4940\ : InMux
    port map (
            O => \N__20714\,
            I => \N__20671\
        );

    \I__4939\ : InMux
    port map (
            O => \N__20713\,
            I => \N__20671\
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__20710\,
            I => bu_rx_data_rdy
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__20707\,
            I => bu_rx_data_rdy
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__20704\,
            I => bu_rx_data_rdy
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__20697\,
            I => bu_rx_data_rdy
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__20692\,
            I => bu_rx_data_rdy
        );

    \I__4933\ : Odrv4
    port map (
            O => \N__20685\,
            I => bu_rx_data_rdy
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__20682\,
            I => bu_rx_data_rdy
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__20679\,
            I => bu_rx_data_rdy
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__20676\,
            I => bu_rx_data_rdy
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__20671\,
            I => bu_rx_data_rdy
        );

    \I__4928\ : CascadeMux
    port map (
            O => \N__20650\,
            I => \Lab_UT.scctrl.N_6_5_cascade_\
        );

    \I__4927\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__20644\,
            I => \Lab_UT.scctrl.N_5_2\
        );

    \I__4925\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20638\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__20638\,
            I => \N__20635\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__20635\,
            I => \Lab_UT.scctrl.N_8_4\
        );

    \I__4922\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20627\
        );

    \I__4921\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20624\
        );

    \I__4920\ : InMux
    port map (
            O => \N__20630\,
            I => \N__20621\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__20627\,
            I => \N__20618\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__20624\,
            I => \N__20615\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__20621\,
            I => \N__20612\
        );

    \I__4916\ : Span4Mux_h
    port map (
            O => \N__20618\,
            I => \N__20608\
        );

    \I__4915\ : Span4Mux_v
    port map (
            O => \N__20615\,
            I => \N__20603\
        );

    \I__4914\ : Span4Mux_v
    port map (
            O => \N__20612\,
            I => \N__20603\
        );

    \I__4913\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20600\
        );

    \I__4912\ : Odrv4
    port map (
            O => \N__20608\,
            I => \Lab_UT.scctrl.N_4ctr\
        );

    \I__4911\ : Odrv4
    port map (
            O => \N__20603\,
            I => \Lab_UT.scctrl.N_4ctr\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__20600\,
            I => \Lab_UT.scctrl.N_4ctr\
        );

    \I__4909\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20590\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__20590\,
            I => \N__20587\
        );

    \I__4907\ : Span4Mux_h
    port map (
            O => \N__20587\,
            I => \N__20584\
        );

    \I__4906\ : Span4Mux_v
    port map (
            O => \N__20584\,
            I => \N__20581\
        );

    \I__4905\ : Odrv4
    port map (
            O => \N__20581\,
            I => \Lab_UT.scctrl.G_23_0_a9_1\
        );

    \I__4904\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20566\
        );

    \I__4903\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20557\
        );

    \I__4902\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20557\
        );

    \I__4901\ : InMux
    port map (
            O => \N__20575\,
            I => \N__20551\
        );

    \I__4900\ : InMux
    port map (
            O => \N__20574\,
            I => \N__20544\
        );

    \I__4899\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20544\
        );

    \I__4898\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20544\
        );

    \I__4897\ : CascadeMux
    port map (
            O => \N__20571\,
            I => \N__20541\
        );

    \I__4896\ : InMux
    port map (
            O => \N__20570\,
            I => \N__20532\
        );

    \I__4895\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20532\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__20566\,
            I => \N__20527\
        );

    \I__4893\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20522\
        );

    \I__4892\ : InMux
    port map (
            O => \N__20564\,
            I => \N__20522\
        );

    \I__4891\ : InMux
    port map (
            O => \N__20563\,
            I => \N__20516\
        );

    \I__4890\ : InMux
    port map (
            O => \N__20562\,
            I => \N__20516\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__20557\,
            I => \N__20513\
        );

    \I__4888\ : InMux
    port map (
            O => \N__20556\,
            I => \N__20505\
        );

    \I__4887\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20505\
        );

    \I__4886\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20505\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20502\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__20544\,
            I => \N__20499\
        );

    \I__4883\ : InMux
    port map (
            O => \N__20541\,
            I => \N__20492\
        );

    \I__4882\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20492\
        );

    \I__4881\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20492\
        );

    \I__4880\ : InMux
    port map (
            O => \N__20538\,
            I => \N__20489\
        );

    \I__4879\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20484\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__20532\,
            I => \N__20481\
        );

    \I__4877\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20478\
        );

    \I__4876\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20475\
        );

    \I__4875\ : Span4Mux_v
    port map (
            O => \N__20527\,
            I => \N__20470\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__20522\,
            I => \N__20470\
        );

    \I__4873\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20467\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__20516\,
            I => \N__20464\
        );

    \I__4871\ : Span12Mux_s10_h
    port map (
            O => \N__20513\,
            I => \N__20459\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__20512\,
            I => \N__20455\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20451\
        );

    \I__4868\ : Span4Mux_s3_h
    port map (
            O => \N__20502\,
            I => \N__20444\
        );

    \I__4867\ : Span4Mux_v
    port map (
            O => \N__20499\,
            I => \N__20444\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__20492\,
            I => \N__20444\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__20489\,
            I => \N__20439\
        );

    \I__4864\ : InMux
    port map (
            O => \N__20488\,
            I => \N__20436\
        );

    \I__4863\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20433\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__20484\,
            I => \N__20418\
        );

    \I__4861\ : Span4Mux_h
    port map (
            O => \N__20481\,
            I => \N__20418\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__20478\,
            I => \N__20418\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__20475\,
            I => \N__20418\
        );

    \I__4858\ : Span4Mux_h
    port map (
            O => \N__20470\,
            I => \N__20418\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__20467\,
            I => \N__20418\
        );

    \I__4856\ : Span4Mux_h
    port map (
            O => \N__20464\,
            I => \N__20418\
        );

    \I__4855\ : InMux
    port map (
            O => \N__20463\,
            I => \N__20415\
        );

    \I__4854\ : InMux
    port map (
            O => \N__20462\,
            I => \N__20412\
        );

    \I__4853\ : Span12Mux_v
    port map (
            O => \N__20459\,
            I => \N__20409\
        );

    \I__4852\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20404\
        );

    \I__4851\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20404\
        );

    \I__4850\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20401\
        );

    \I__4849\ : Span4Mux_s3_h
    port map (
            O => \N__20451\,
            I => \N__20396\
        );

    \I__4848\ : Span4Mux_v
    port map (
            O => \N__20444\,
            I => \N__20396\
        );

    \I__4847\ : InMux
    port map (
            O => \N__20443\,
            I => \N__20391\
        );

    \I__4846\ : InMux
    port map (
            O => \N__20442\,
            I => \N__20391\
        );

    \I__4845\ : Span12Mux_s2_v
    port map (
            O => \N__20439\,
            I => \N__20382\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__20436\,
            I => \N__20382\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__20433\,
            I => \N__20382\
        );

    \I__4842\ : Sp12to4
    port map (
            O => \N__20418\,
            I => \N__20382\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__20415\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__20412\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__4839\ : Odrv12
    port map (
            O => \N__20409\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__20404\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__20401\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__20396\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__20391\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__4834\ : Odrv12
    port map (
            O => \N__20382\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__4833\ : InMux
    port map (
            O => \N__20365\,
            I => \N__20356\
        );

    \I__4832\ : InMux
    port map (
            O => \N__20364\,
            I => \N__20356\
        );

    \I__4831\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20356\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__20356\,
            I => \N__20353\
        );

    \I__4829\ : Odrv4
    port map (
            O => \N__20353\,
            I => \Lab_UT.scctrl.g0_i_a8_4_1\
        );

    \I__4828\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20345\
        );

    \I__4827\ : CascadeMux
    port map (
            O => \N__20349\,
            I => \N__20342\
        );

    \I__4826\ : InMux
    port map (
            O => \N__20348\,
            I => \N__20338\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__20345\,
            I => \N__20335\
        );

    \I__4824\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20332\
        );

    \I__4823\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20328\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__20338\,
            I => \N__20325\
        );

    \I__4821\ : Span4Mux_s2_h
    port map (
            O => \N__20335\,
            I => \N__20320\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__20332\,
            I => \N__20320\
        );

    \I__4819\ : InMux
    port map (
            O => \N__20331\,
            I => \N__20317\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__20328\,
            I => \N__20312\
        );

    \I__4817\ : Span4Mux_h
    port map (
            O => \N__20325\,
            I => \N__20312\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__20320\,
            I => \N__20309\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20303\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__20312\,
            I => \N__20303\
        );

    \I__4813\ : Span4Mux_v
    port map (
            O => \N__20309\,
            I => \N__20300\
        );

    \I__4812\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20297\
        );

    \I__4811\ : Span4Mux_v
    port map (
            O => \N__20303\,
            I => \N__20294\
        );

    \I__4810\ : Span4Mux_v
    port map (
            O => \N__20300\,
            I => \N__20291\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__20297\,
            I => \Lab_UT.scctrl.next_state_0_2\
        );

    \I__4808\ : Odrv4
    port map (
            O => \N__20294\,
            I => \Lab_UT.scctrl.next_state_0_2\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__20291\,
            I => \Lab_UT.scctrl.next_state_0_2\
        );

    \I__4806\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20279\
        );

    \I__4805\ : InMux
    port map (
            O => \N__20283\,
            I => \N__20276\
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__20282\,
            I => \N__20273\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__20279\,
            I => \N__20264\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__20276\,
            I => \N__20261\
        );

    \I__4801\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20258\
        );

    \I__4800\ : CascadeMux
    port map (
            O => \N__20272\,
            I => \N__20253\
        );

    \I__4799\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20250\
        );

    \I__4798\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20247\
        );

    \I__4797\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20244\
        );

    \I__4796\ : InMux
    port map (
            O => \N__20268\,
            I => \N__20240\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20237\
        );

    \I__4794\ : Span4Mux_v
    port map (
            O => \N__20264\,
            I => \N__20230\
        );

    \I__4793\ : Span4Mux_h
    port map (
            O => \N__20261\,
            I => \N__20230\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__20258\,
            I => \N__20230\
        );

    \I__4791\ : CascadeMux
    port map (
            O => \N__20257\,
            I => \N__20226\
        );

    \I__4790\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20223\
        );

    \I__4789\ : InMux
    port map (
            O => \N__20253\,
            I => \N__20219\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__20250\,
            I => \N__20216\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__20247\,
            I => \N__20213\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__20244\,
            I => \N__20210\
        );

    \I__4785\ : InMux
    port map (
            O => \N__20243\,
            I => \N__20206\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__20240\,
            I => \N__20201\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__20237\,
            I => \N__20201\
        );

    \I__4782\ : Span4Mux_v
    port map (
            O => \N__20230\,
            I => \N__20198\
        );

    \I__4781\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20195\
        );

    \I__4780\ : InMux
    port map (
            O => \N__20226\,
            I => \N__20192\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__20223\,
            I => \N__20189\
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__20222\,
            I => \N__20185\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__20219\,
            I => \N__20179\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__20216\,
            I => \N__20179\
        );

    \I__4775\ : Span4Mux_v
    port map (
            O => \N__20213\,
            I => \N__20174\
        );

    \I__4774\ : Span4Mux_s1_h
    port map (
            O => \N__20210\,
            I => \N__20174\
        );

    \I__4773\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20171\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__20206\,
            I => \N__20168\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__20201\,
            I => \N__20165\
        );

    \I__4770\ : Span4Mux_h
    port map (
            O => \N__20198\,
            I => \N__20156\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__20195\,
            I => \N__20156\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__20192\,
            I => \N__20156\
        );

    \I__4767\ : Span4Mux_s3_v
    port map (
            O => \N__20189\,
            I => \N__20152\
        );

    \I__4766\ : InMux
    port map (
            O => \N__20188\,
            I => \N__20147\
        );

    \I__4765\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20147\
        );

    \I__4764\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20144\
        );

    \I__4763\ : Span4Mux_h
    port map (
            O => \N__20179\,
            I => \N__20137\
        );

    \I__4762\ : Span4Mux_h
    port map (
            O => \N__20174\,
            I => \N__20137\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__20171\,
            I => \N__20137\
        );

    \I__4760\ : Span4Mux_h
    port map (
            O => \N__20168\,
            I => \N__20132\
        );

    \I__4759\ : Span4Mux_v
    port map (
            O => \N__20165\,
            I => \N__20132\
        );

    \I__4758\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20127\
        );

    \I__4757\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20127\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__20156\,
            I => \N__20124\
        );

    \I__4755\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20121\
        );

    \I__4754\ : Sp12to4
    port map (
            O => \N__20152\,
            I => \N__20116\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__20147\,
            I => \N__20116\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__20144\,
            I => \N__20111\
        );

    \I__4751\ : Span4Mux_v
    port map (
            O => \N__20137\,
            I => \N__20111\
        );

    \I__4750\ : Odrv4
    port map (
            O => \N__20132\,
            I => rst_i_3
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__20127\,
            I => rst_i_3
        );

    \I__4748\ : Odrv4
    port map (
            O => \N__20124\,
            I => rst_i_3
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__20121\,
            I => rst_i_3
        );

    \I__4746\ : Odrv12
    port map (
            O => \N__20116\,
            I => rst_i_3
        );

    \I__4745\ : Odrv4
    port map (
            O => \N__20111\,
            I => rst_i_3
        );

    \I__4744\ : InMux
    port map (
            O => \N__20098\,
            I => \N__20085\
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__20097\,
            I => \N__20072\
        );

    \I__4742\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20066\
        );

    \I__4741\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20063\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__20094\,
            I => \N__20056\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__20093\,
            I => \N__20053\
        );

    \I__4738\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20041\
        );

    \I__4737\ : InMux
    port map (
            O => \N__20091\,
            I => \N__20041\
        );

    \I__4736\ : InMux
    port map (
            O => \N__20090\,
            I => \N__20041\
        );

    \I__4735\ : InMux
    port map (
            O => \N__20089\,
            I => \N__20041\
        );

    \I__4734\ : InMux
    port map (
            O => \N__20088\,
            I => \N__20038\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__20085\,
            I => \N__20035\
        );

    \I__4732\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20028\
        );

    \I__4731\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20028\
        );

    \I__4730\ : InMux
    port map (
            O => \N__20082\,
            I => \N__20028\
        );

    \I__4729\ : InMux
    port map (
            O => \N__20081\,
            I => \N__20021\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20080\,
            I => \N__20021\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20021\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20078\,
            I => \N__20015\
        );

    \I__4725\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20012\
        );

    \I__4724\ : InMux
    port map (
            O => \N__20076\,
            I => \N__20009\
        );

    \I__4723\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20002\
        );

    \I__4722\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20002\
        );

    \I__4721\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20002\
        );

    \I__4720\ : InMux
    port map (
            O => \N__20070\,
            I => \N__19999\
        );

    \I__4719\ : CascadeMux
    port map (
            O => \N__20069\,
            I => \N__19993\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__20066\,
            I => \N__19987\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__20063\,
            I => \N__19987\
        );

    \I__4716\ : InMux
    port map (
            O => \N__20062\,
            I => \N__19984\
        );

    \I__4715\ : InMux
    port map (
            O => \N__20061\,
            I => \N__19981\
        );

    \I__4714\ : InMux
    port map (
            O => \N__20060\,
            I => \N__19978\
        );

    \I__4713\ : InMux
    port map (
            O => \N__20059\,
            I => \N__19973\
        );

    \I__4712\ : InMux
    port map (
            O => \N__20056\,
            I => \N__19973\
        );

    \I__4711\ : InMux
    port map (
            O => \N__20053\,
            I => \N__19958\
        );

    \I__4710\ : InMux
    port map (
            O => \N__20052\,
            I => \N__19955\
        );

    \I__4709\ : InMux
    port map (
            O => \N__20051\,
            I => \N__19952\
        );

    \I__4708\ : InMux
    port map (
            O => \N__20050\,
            I => \N__19949\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__20041\,
            I => \N__19944\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__20038\,
            I => \N__19944\
        );

    \I__4705\ : Span4Mux_v
    port map (
            O => \N__20035\,
            I => \N__19941\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__20028\,
            I => \N__19936\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__20021\,
            I => \N__19936\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20020\,
            I => \N__19931\
        );

    \I__4701\ : InMux
    port map (
            O => \N__20019\,
            I => \N__19931\
        );

    \I__4700\ : InMux
    port map (
            O => \N__20018\,
            I => \N__19928\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__20015\,
            I => \N__19923\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__20012\,
            I => \N__19923\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__20009\,
            I => \N__19918\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__20002\,
            I => \N__19918\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__19999\,
            I => \N__19912\
        );

    \I__4694\ : InMux
    port map (
            O => \N__19998\,
            I => \N__19909\
        );

    \I__4693\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19904\
        );

    \I__4692\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19904\
        );

    \I__4691\ : InMux
    port map (
            O => \N__19993\,
            I => \N__19899\
        );

    \I__4690\ : InMux
    port map (
            O => \N__19992\,
            I => \N__19899\
        );

    \I__4689\ : Span4Mux_v
    port map (
            O => \N__19987\,
            I => \N__19894\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__19984\,
            I => \N__19894\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__19981\,
            I => \N__19889\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__19978\,
            I => \N__19889\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__19973\,
            I => \N__19886\
        );

    \I__4684\ : InMux
    port map (
            O => \N__19972\,
            I => \N__19881\
        );

    \I__4683\ : InMux
    port map (
            O => \N__19971\,
            I => \N__19881\
        );

    \I__4682\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19872\
        );

    \I__4681\ : InMux
    port map (
            O => \N__19969\,
            I => \N__19869\
        );

    \I__4680\ : InMux
    port map (
            O => \N__19968\,
            I => \N__19866\
        );

    \I__4679\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19857\
        );

    \I__4678\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19857\
        );

    \I__4677\ : InMux
    port map (
            O => \N__19965\,
            I => \N__19857\
        );

    \I__4676\ : InMux
    port map (
            O => \N__19964\,
            I => \N__19857\
        );

    \I__4675\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19850\
        );

    \I__4674\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19850\
        );

    \I__4673\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19850\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__19958\,
            I => \N__19847\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__19955\,
            I => \N__19836\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19836\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__19949\,
            I => \N__19836\
        );

    \I__4668\ : Span4Mux_v
    port map (
            O => \N__19944\,
            I => \N__19836\
        );

    \I__4667\ : Span4Mux_h
    port map (
            O => \N__19941\,
            I => \N__19836\
        );

    \I__4666\ : Span4Mux_h
    port map (
            O => \N__19936\,
            I => \N__19831\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__19931\,
            I => \N__19828\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__19928\,
            I => \N__19821\
        );

    \I__4663\ : Span4Mux_v
    port map (
            O => \N__19923\,
            I => \N__19821\
        );

    \I__4662\ : Span4Mux_v
    port map (
            O => \N__19918\,
            I => \N__19821\
        );

    \I__4661\ : InMux
    port map (
            O => \N__19917\,
            I => \N__19814\
        );

    \I__4660\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19814\
        );

    \I__4659\ : InMux
    port map (
            O => \N__19915\,
            I => \N__19814\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__19912\,
            I => \N__19807\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__19909\,
            I => \N__19807\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__19904\,
            I => \N__19807\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__19899\,
            I => \N__19804\
        );

    \I__4654\ : Span4Mux_h
    port map (
            O => \N__19894\,
            I => \N__19801\
        );

    \I__4653\ : Span4Mux_h
    port map (
            O => \N__19889\,
            I => \N__19796\
        );

    \I__4652\ : Span4Mux_v
    port map (
            O => \N__19886\,
            I => \N__19796\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__19881\,
            I => \N__19793\
        );

    \I__4650\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19788\
        );

    \I__4649\ : InMux
    port map (
            O => \N__19879\,
            I => \N__19788\
        );

    \I__4648\ : InMux
    port map (
            O => \N__19878\,
            I => \N__19781\
        );

    \I__4647\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19781\
        );

    \I__4646\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19781\
        );

    \I__4645\ : InMux
    port map (
            O => \N__19875\,
            I => \N__19778\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__19872\,
            I => \N__19775\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__19869\,
            I => \N__19762\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__19866\,
            I => \N__19762\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19762\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__19850\,
            I => \N__19762\
        );

    \I__4639\ : Span4Mux_v
    port map (
            O => \N__19847\,
            I => \N__19762\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__19836\,
            I => \N__19762\
        );

    \I__4637\ : InMux
    port map (
            O => \N__19835\,
            I => \N__19757\
        );

    \I__4636\ : InMux
    port map (
            O => \N__19834\,
            I => \N__19757\
        );

    \I__4635\ : Span4Mux_v
    port map (
            O => \N__19831\,
            I => \N__19752\
        );

    \I__4634\ : Span4Mux_s2_h
    port map (
            O => \N__19828\,
            I => \N__19752\
        );

    \I__4633\ : Span4Mux_v
    port map (
            O => \N__19821\,
            I => \N__19743\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__19814\,
            I => \N__19743\
        );

    \I__4631\ : Span4Mux_v
    port map (
            O => \N__19807\,
            I => \N__19743\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__19804\,
            I => \N__19743\
        );

    \I__4629\ : Span4Mux_v
    port map (
            O => \N__19801\,
            I => \N__19736\
        );

    \I__4628\ : Span4Mux_v
    port map (
            O => \N__19796\,
            I => \N__19736\
        );

    \I__4627\ : Span4Mux_s2_h
    port map (
            O => \N__19793\,
            I => \N__19736\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__19788\,
            I => \Lab_UT_scctrl_N_221_0\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__19781\,
            I => \Lab_UT_scctrl_N_221_0\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__19778\,
            I => \Lab_UT_scctrl_N_221_0\
        );

    \I__4623\ : Odrv12
    port map (
            O => \N__19775\,
            I => \Lab_UT_scctrl_N_221_0\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__19762\,
            I => \Lab_UT_scctrl_N_221_0\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__19757\,
            I => \Lab_UT_scctrl_N_221_0\
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__19752\,
            I => \Lab_UT_scctrl_N_221_0\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__19743\,
            I => \Lab_UT_scctrl_N_221_0\
        );

    \I__4618\ : Odrv4
    port map (
            O => \N__19736\,
            I => \Lab_UT_scctrl_N_221_0\
        );

    \I__4617\ : InMux
    port map (
            O => \N__19717\,
            I => \N__19711\
        );

    \I__4616\ : InMux
    port map (
            O => \N__19716\,
            I => \N__19711\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__19711\,
            I => \N__19708\
        );

    \I__4614\ : Odrv12
    port map (
            O => \N__19708\,
            I => \Lab_UT.scctrl.G_21_i_0\
        );

    \I__4613\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19700\
        );

    \I__4612\ : CascadeMux
    port map (
            O => \N__19704\,
            I => \N__19692\
        );

    \I__4611\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19688\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__19700\,
            I => \N__19685\
        );

    \I__4609\ : InMux
    port map (
            O => \N__19699\,
            I => \N__19680\
        );

    \I__4608\ : InMux
    port map (
            O => \N__19698\,
            I => \N__19680\
        );

    \I__4607\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19675\
        );

    \I__4606\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19670\
        );

    \I__4605\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19670\
        );

    \I__4604\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19667\
        );

    \I__4603\ : CascadeMux
    port map (
            O => \N__19691\,
            I => \N__19663\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__19688\,
            I => \N__19659\
        );

    \I__4601\ : Span4Mux_v
    port map (
            O => \N__19685\,
            I => \N__19655\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__19680\,
            I => \N__19651\
        );

    \I__4599\ : InMux
    port map (
            O => \N__19679\,
            I => \N__19646\
        );

    \I__4598\ : InMux
    port map (
            O => \N__19678\,
            I => \N__19646\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__19675\,
            I => \N__19643\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__19670\,
            I => \N__19640\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__19667\,
            I => \N__19637\
        );

    \I__4594\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19632\
        );

    \I__4593\ : InMux
    port map (
            O => \N__19663\,
            I => \N__19632\
        );

    \I__4592\ : InMux
    port map (
            O => \N__19662\,
            I => \N__19629\
        );

    \I__4591\ : Span4Mux_h
    port map (
            O => \N__19659\,
            I => \N__19625\
        );

    \I__4590\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19622\
        );

    \I__4589\ : IoSpan4Mux
    port map (
            O => \N__19655\,
            I => \N__19618\
        );

    \I__4588\ : InMux
    port map (
            O => \N__19654\,
            I => \N__19615\
        );

    \I__4587\ : Span4Mux_s3_v
    port map (
            O => \N__19651\,
            I => \N__19612\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19605\
        );

    \I__4585\ : Span4Mux_h
    port map (
            O => \N__19643\,
            I => \N__19605\
        );

    \I__4584\ : Span4Mux_v
    port map (
            O => \N__19640\,
            I => \N__19605\
        );

    \I__4583\ : Span4Mux_s2_v
    port map (
            O => \N__19637\,
            I => \N__19598\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__19632\,
            I => \N__19598\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__19629\,
            I => \N__19598\
        );

    \I__4580\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19595\
        );

    \I__4579\ : Span4Mux_v
    port map (
            O => \N__19625\,
            I => \N__19592\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__19622\,
            I => \N__19589\
        );

    \I__4577\ : InMux
    port map (
            O => \N__19621\,
            I => \N__19586\
        );

    \I__4576\ : Span4Mux_s1_h
    port map (
            O => \N__19618\,
            I => \N__19579\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__19615\,
            I => \N__19579\
        );

    \I__4574\ : Span4Mux_h
    port map (
            O => \N__19612\,
            I => \N__19579\
        );

    \I__4573\ : Span4Mux_v
    port map (
            O => \N__19605\,
            I => \N__19574\
        );

    \I__4572\ : Span4Mux_v
    port map (
            O => \N__19598\,
            I => \N__19574\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__19595\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__19592\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4569\ : Odrv4
    port map (
            O => \N__19589\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__19586\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4567\ : Odrv4
    port map (
            O => \N__19579\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__19574\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4565\ : CascadeMux
    port map (
            O => \N__19561\,
            I => \N__19557\
        );

    \I__4564\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19547\
        );

    \I__4563\ : InMux
    port map (
            O => \N__19557\,
            I => \N__19544\
        );

    \I__4562\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19539\
        );

    \I__4561\ : InMux
    port map (
            O => \N__19555\,
            I => \N__19539\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__19554\,
            I => \N__19534\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__19553\,
            I => \N__19531\
        );

    \I__4558\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19525\
        );

    \I__4557\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19525\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__19550\,
            I => \N__19522\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__19547\,
            I => \N__19518\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__19544\,
            I => \N__19515\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__19539\,
            I => \N__19512\
        );

    \I__4552\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19509\
        );

    \I__4551\ : InMux
    port map (
            O => \N__19537\,
            I => \N__19506\
        );

    \I__4550\ : InMux
    port map (
            O => \N__19534\,
            I => \N__19503\
        );

    \I__4549\ : InMux
    port map (
            O => \N__19531\,
            I => \N__19500\
        );

    \I__4548\ : InMux
    port map (
            O => \N__19530\,
            I => \N__19497\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__19525\,
            I => \N__19494\
        );

    \I__4546\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19491\
        );

    \I__4545\ : InMux
    port map (
            O => \N__19521\,
            I => \N__19488\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__19518\,
            I => \N__19474\
        );

    \I__4543\ : Span4Mux_h
    port map (
            O => \N__19515\,
            I => \N__19474\
        );

    \I__4542\ : Span4Mux_v
    port map (
            O => \N__19512\,
            I => \N__19474\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__19509\,
            I => \N__19474\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__19506\,
            I => \N__19474\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__19503\,
            I => \N__19471\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__19500\,
            I => \N__19468\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__19497\,
            I => \N__19463\
        );

    \I__4536\ : Span4Mux_h
    port map (
            O => \N__19494\,
            I => \N__19463\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__19491\,
            I => \N__19460\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__19488\,
            I => \N__19457\
        );

    \I__4533\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19450\
        );

    \I__4532\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19450\
        );

    \I__4531\ : InMux
    port map (
            O => \N__19485\,
            I => \N__19450\
        );

    \I__4530\ : Span4Mux_h
    port map (
            O => \N__19474\,
            I => \N__19447\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__19471\,
            I => \N__19440\
        );

    \I__4528\ : Span4Mux_h
    port map (
            O => \N__19468\,
            I => \N__19440\
        );

    \I__4527\ : Span4Mux_v
    port map (
            O => \N__19463\,
            I => \N__19440\
        );

    \I__4526\ : Odrv4
    port map (
            O => \N__19460\,
            I => \Lab_UT.state_2\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__19457\,
            I => \Lab_UT.state_2\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__19450\,
            I => \Lab_UT.state_2\
        );

    \I__4523\ : Odrv4
    port map (
            O => \N__19447\,
            I => \Lab_UT.state_2\
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__19440\,
            I => \Lab_UT.state_2\
        );

    \I__4521\ : InMux
    port map (
            O => \N__19429\,
            I => \N__19426\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__19426\,
            I => \N__19422\
        );

    \I__4519\ : InMux
    port map (
            O => \N__19425\,
            I => \N__19419\
        );

    \I__4518\ : Span4Mux_s2_h
    port map (
            O => \N__19422\,
            I => \N__19416\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__19419\,
            I => \N__19413\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__19416\,
            I => \Lab_UT.scctrl.N_11_1\
        );

    \I__4515\ : Odrv4
    port map (
            O => \N__19413\,
            I => \Lab_UT.scctrl.N_11_1\
        );

    \I__4514\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19405\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__19405\,
            I => \N__19402\
        );

    \I__4512\ : Span4Mux_s3_h
    port map (
            O => \N__19402\,
            I => \N__19399\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__19399\,
            I => \Lab_UT.scctrl.N_12_2\
        );

    \I__4510\ : CascadeMux
    port map (
            O => \N__19396\,
            I => \Lab_UT.scctrl.G_24_i_a4_1_cascade_\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__19393\,
            I => \N__19390\
        );

    \I__4508\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19387\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__19387\,
            I => \N__19384\
        );

    \I__4506\ : Odrv4
    port map (
            O => \N__19384\,
            I => \Lab_UT.scctrl.G_21_i_a7_0_1\
        );

    \I__4505\ : InMux
    port map (
            O => \N__19381\,
            I => \N__19372\
        );

    \I__4504\ : InMux
    port map (
            O => \N__19380\,
            I => \N__19372\
        );

    \I__4503\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19372\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__19372\,
            I => \N__19368\
        );

    \I__4501\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19365\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__19368\,
            I => \Lab_UT.scctrl.N_9_2\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__19365\,
            I => \Lab_UT.scctrl.N_9_2\
        );

    \I__4498\ : CascadeMux
    port map (
            O => \N__19360\,
            I => \N__19356\
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__19359\,
            I => \N__19353\
        );

    \I__4496\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19348\
        );

    \I__4495\ : InMux
    port map (
            O => \N__19353\,
            I => \N__19348\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__19348\,
            I => \Lab_UT.scctrl.G_21_i_2\
        );

    \I__4493\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19335\
        );

    \I__4492\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19335\
        );

    \I__4491\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19335\
        );

    \I__4490\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19332\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__19335\,
            I => \Lab_UT.scctrl.N_8_2\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__19332\,
            I => \Lab_UT.scctrl.N_8_2\
        );

    \I__4487\ : CascadeMux
    port map (
            O => \N__19327\,
            I => \N__19324\
        );

    \I__4486\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19320\
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__19323\,
            I => \N__19316\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__19320\,
            I => \N__19311\
        );

    \I__4483\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19306\
        );

    \I__4482\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19303\
        );

    \I__4481\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19300\
        );

    \I__4480\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19297\
        );

    \I__4479\ : Span4Mux_s2_h
    port map (
            O => \N__19311\,
            I => \N__19294\
        );

    \I__4478\ : InMux
    port map (
            O => \N__19310\,
            I => \N__19289\
        );

    \I__4477\ : InMux
    port map (
            O => \N__19309\,
            I => \N__19286\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__19306\,
            I => \N__19281\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__19303\,
            I => \N__19281\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__19300\,
            I => \N__19278\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__19297\,
            I => \N__19275\
        );

    \I__4472\ : Span4Mux_v
    port map (
            O => \N__19294\,
            I => \N__19272\
        );

    \I__4471\ : InMux
    port map (
            O => \N__19293\,
            I => \N__19269\
        );

    \I__4470\ : InMux
    port map (
            O => \N__19292\,
            I => \N__19266\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__19289\,
            I => \N__19263\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__19286\,
            I => \N__19254\
        );

    \I__4467\ : Span4Mux_s3_h
    port map (
            O => \N__19281\,
            I => \N__19254\
        );

    \I__4466\ : Span4Mux_v
    port map (
            O => \N__19278\,
            I => \N__19254\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__19275\,
            I => \N__19254\
        );

    \I__4464\ : Odrv4
    port map (
            O => \N__19272\,
            I => \Lab_UT.state_i_3_0_rep1\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__19269\,
            I => \Lab_UT.state_i_3_0_rep1\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__19266\,
            I => \Lab_UT.state_i_3_0_rep1\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__19263\,
            I => \Lab_UT.state_i_3_0_rep1\
        );

    \I__4460\ : Odrv4
    port map (
            O => \N__19254\,
            I => \Lab_UT.state_i_3_0_rep1\
        );

    \I__4459\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19240\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__19240\,
            I => \N__19234\
        );

    \I__4457\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19231\
        );

    \I__4456\ : InMux
    port map (
            O => \N__19238\,
            I => \N__19228\
        );

    \I__4455\ : InMux
    port map (
            O => \N__19237\,
            I => \N__19225\
        );

    \I__4454\ : Span4Mux_v
    port map (
            O => \N__19234\,
            I => \N__19220\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__19231\,
            I => \N__19220\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__19228\,
            I => \N__19216\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__19225\,
            I => \N__19213\
        );

    \I__4450\ : Span4Mux_h
    port map (
            O => \N__19220\,
            I => \N__19207\
        );

    \I__4449\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19204\
        );

    \I__4448\ : Span12Mux_s4_h
    port map (
            O => \N__19216\,
            I => \N__19199\
        );

    \I__4447\ : Span12Mux_s5_v
    port map (
            O => \N__19213\,
            I => \N__19199\
        );

    \I__4446\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19194\
        );

    \I__4445\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19194\
        );

    \I__4444\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19191\
        );

    \I__4443\ : Odrv4
    port map (
            O => \N__19207\,
            I => \Lab_UT.state_i_3_2_rep1\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__19204\,
            I => \Lab_UT.state_i_3_2_rep1\
        );

    \I__4441\ : Odrv12
    port map (
            O => \N__19199\,
            I => \Lab_UT.state_i_3_2_rep1\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__19194\,
            I => \Lab_UT.state_i_3_2_rep1\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__19191\,
            I => \Lab_UT.state_i_3_2_rep1\
        );

    \I__4438\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19177\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__19177\,
            I => \N__19174\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__19174\,
            I => \Lab_UT.scctrl.g0_1_4_1\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__19171\,
            I => \Lab_UT.scctrl.g0_i_a7_0_1_cascade_\
        );

    \I__4434\ : InMux
    port map (
            O => \N__19168\,
            I => \N__19158\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__19167\,
            I => \N__19152\
        );

    \I__4432\ : InMux
    port map (
            O => \N__19166\,
            I => \N__19144\
        );

    \I__4431\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19139\
        );

    \I__4430\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19139\
        );

    \I__4429\ : InMux
    port map (
            O => \N__19163\,
            I => \N__19134\
        );

    \I__4428\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19134\
        );

    \I__4427\ : InMux
    port map (
            O => \N__19161\,
            I => \N__19131\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__19158\,
            I => \N__19128\
        );

    \I__4425\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19125\
        );

    \I__4424\ : InMux
    port map (
            O => \N__19156\,
            I => \N__19122\
        );

    \I__4423\ : InMux
    port map (
            O => \N__19155\,
            I => \N__19119\
        );

    \I__4422\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19113\
        );

    \I__4421\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19113\
        );

    \I__4420\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19110\
        );

    \I__4419\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19102\
        );

    \I__4418\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19102\
        );

    \I__4417\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19098\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__19144\,
            I => \N__19091\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__19139\,
            I => \N__19091\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__19134\,
            I => \N__19087\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__19131\,
            I => \N__19084\
        );

    \I__4412\ : Span4Mux_v
    port map (
            O => \N__19128\,
            I => \N__19079\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__19125\,
            I => \N__19079\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__19122\,
            I => \N__19076\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__19119\,
            I => \N__19073\
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__19118\,
            I => \N__19070\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__19113\,
            I => \N__19066\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__19110\,
            I => \N__19063\
        );

    \I__4405\ : InMux
    port map (
            O => \N__19109\,
            I => \N__19058\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19108\,
            I => \N__19058\
        );

    \I__4403\ : InMux
    port map (
            O => \N__19107\,
            I => \N__19055\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__19102\,
            I => \N__19052\
        );

    \I__4401\ : InMux
    port map (
            O => \N__19101\,
            I => \N__19049\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__19098\,
            I => \N__19046\
        );

    \I__4399\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19041\
        );

    \I__4398\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19041\
        );

    \I__4397\ : Span4Mux_h
    port map (
            O => \N__19091\,
            I => \N__19038\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19090\,
            I => \N__19035\
        );

    \I__4395\ : Span4Mux_v
    port map (
            O => \N__19087\,
            I => \N__19032\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__19084\,
            I => \N__19027\
        );

    \I__4393\ : Span4Mux_h
    port map (
            O => \N__19079\,
            I => \N__19027\
        );

    \I__4392\ : Span4Mux_v
    port map (
            O => \N__19076\,
            I => \N__19022\
        );

    \I__4391\ : Span4Mux_s1_h
    port map (
            O => \N__19073\,
            I => \N__19022\
        );

    \I__4390\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19017\
        );

    \I__4389\ : InMux
    port map (
            O => \N__19069\,
            I => \N__19017\
        );

    \I__4388\ : Span12Mux_s5_h
    port map (
            O => \N__19066\,
            I => \N__19010\
        );

    \I__4387\ : Sp12to4
    port map (
            O => \N__19063\,
            I => \N__19010\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__19058\,
            I => \N__19010\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__19055\,
            I => \N__19003\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__19052\,
            I => \N__19003\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__19049\,
            I => \N__19003\
        );

    \I__4382\ : Odrv4
    port map (
            O => \N__19046\,
            I => \Lab_UT.de_hex_0\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__19041\,
            I => \Lab_UT.de_hex_0\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__19038\,
            I => \Lab_UT.de_hex_0\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__19035\,
            I => \Lab_UT.de_hex_0\
        );

    \I__4378\ : Odrv4
    port map (
            O => \N__19032\,
            I => \Lab_UT.de_hex_0\
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__19027\,
            I => \Lab_UT.de_hex_0\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__19022\,
            I => \Lab_UT.de_hex_0\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__19017\,
            I => \Lab_UT.de_hex_0\
        );

    \I__4374\ : Odrv12
    port map (
            O => \N__19010\,
            I => \Lab_UT.de_hex_0\
        );

    \I__4373\ : Odrv4
    port map (
            O => \N__19003\,
            I => \Lab_UT.de_hex_0\
        );

    \I__4372\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18979\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__18979\,
            I => \N__18976\
        );

    \I__4370\ : Odrv12
    port map (
            O => \N__18976\,
            I => \Lab_UT.scctrl.N_10_0\
        );

    \I__4369\ : CascadeMux
    port map (
            O => \N__18973\,
            I => \Lab_UT.scctrl.g0_7_a13_1_1_cascade_\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__18970\,
            I => \Lab_UT.scctrl.N_7_cascade_\
        );

    \I__4367\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18964\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__18964\,
            I => \N__18961\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__18961\,
            I => \N__18958\
        );

    \I__4364\ : Odrv4
    port map (
            O => \N__18958\,
            I => \Lab_UT.scctrl.g0_6\
        );

    \I__4363\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18948\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__18954\,
            I => \N__18943\
        );

    \I__4361\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18940\
        );

    \I__4360\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18935\
        );

    \I__4359\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18932\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__18948\,
            I => \N__18929\
        );

    \I__4357\ : InMux
    port map (
            O => \N__18947\,
            I => \N__18926\
        );

    \I__4356\ : InMux
    port map (
            O => \N__18946\,
            I => \N__18923\
        );

    \I__4355\ : InMux
    port map (
            O => \N__18943\,
            I => \N__18919\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__18940\,
            I => \N__18915\
        );

    \I__4353\ : InMux
    port map (
            O => \N__18939\,
            I => \N__18910\
        );

    \I__4352\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18907\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__18935\,
            I => \N__18904\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__18932\,
            I => \N__18899\
        );

    \I__4349\ : Span4Mux_s3_v
    port map (
            O => \N__18929\,
            I => \N__18899\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__18926\,
            I => \N__18896\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__18923\,
            I => \N__18893\
        );

    \I__4346\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18890\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__18919\,
            I => \N__18887\
        );

    \I__4344\ : InMux
    port map (
            O => \N__18918\,
            I => \N__18884\
        );

    \I__4343\ : Span4Mux_s2_v
    port map (
            O => \N__18915\,
            I => \N__18881\
        );

    \I__4342\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18876\
        );

    \I__4341\ : InMux
    port map (
            O => \N__18913\,
            I => \N__18876\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__18910\,
            I => \N__18873\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__18907\,
            I => \N__18870\
        );

    \I__4338\ : Span4Mux_h
    port map (
            O => \N__18904\,
            I => \N__18864\
        );

    \I__4337\ : Span4Mux_h
    port map (
            O => \N__18899\,
            I => \N__18864\
        );

    \I__4336\ : Span4Mux_v
    port map (
            O => \N__18896\,
            I => \N__18859\
        );

    \I__4335\ : Span4Mux_h
    port map (
            O => \N__18893\,
            I => \N__18859\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__18890\,
            I => \N__18855\
        );

    \I__4333\ : Span4Mux_v
    port map (
            O => \N__18887\,
            I => \N__18844\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__18884\,
            I => \N__18844\
        );

    \I__4331\ : Span4Mux_v
    port map (
            O => \N__18881\,
            I => \N__18844\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__18876\,
            I => \N__18844\
        );

    \I__4329\ : Span4Mux_v
    port map (
            O => \N__18873\,
            I => \N__18844\
        );

    \I__4328\ : Span4Mux_s2_v
    port map (
            O => \N__18870\,
            I => \N__18841\
        );

    \I__4327\ : InMux
    port map (
            O => \N__18869\,
            I => \N__18838\
        );

    \I__4326\ : Span4Mux_v
    port map (
            O => \N__18864\,
            I => \N__18833\
        );

    \I__4325\ : Span4Mux_h
    port map (
            O => \N__18859\,
            I => \N__18833\
        );

    \I__4324\ : InMux
    port map (
            O => \N__18858\,
            I => \N__18830\
        );

    \I__4323\ : Span4Mux_v
    port map (
            O => \N__18855\,
            I => \N__18823\
        );

    \I__4322\ : Span4Mux_h
    port map (
            O => \N__18844\,
            I => \N__18823\
        );

    \I__4321\ : Span4Mux_v
    port map (
            O => \N__18841\,
            I => \N__18823\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__18838\,
            I => rst
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__18833\,
            I => rst
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__18830\,
            I => rst
        );

    \I__4317\ : Odrv4
    port map (
            O => \N__18823\,
            I => rst
        );

    \I__4316\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18811\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__18811\,
            I => \N__18808\
        );

    \I__4314\ : Odrv12
    port map (
            O => \N__18808\,
            I => \Lab_UT.scctrl.g1_i_a7_2Z0Z_3\
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__18805\,
            I => \Lab_UT.scctrl.N_10_1_cascade_\
        );

    \I__4312\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18799\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__18799\,
            I => \N__18796\
        );

    \I__4310\ : Span4Mux_v
    port map (
            O => \N__18796\,
            I => \N__18793\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__18793\,
            I => \Lab_UT.scctrl.g1_i_2\
        );

    \I__4308\ : InMux
    port map (
            O => \N__18790\,
            I => \N__18787\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__18787\,
            I => \Lab_UT.scctrl.N_7_4\
        );

    \I__4306\ : InMux
    port map (
            O => \N__18784\,
            I => \N__18777\
        );

    \I__4305\ : InMux
    port map (
            O => \N__18783\,
            I => \N__18774\
        );

    \I__4304\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18766\
        );

    \I__4303\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18766\
        );

    \I__4302\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18760\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__18777\,
            I => \N__18755\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__18774\,
            I => \N__18755\
        );

    \I__4299\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18752\
        );

    \I__4298\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18745\
        );

    \I__4297\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18742\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__18766\,
            I => \N__18739\
        );

    \I__4295\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18736\
        );

    \I__4294\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18731\
        );

    \I__4293\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18731\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__18760\,
            I => \N__18725\
        );

    \I__4291\ : Span4Mux_s3_h
    port map (
            O => \N__18755\,
            I => \N__18722\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__18752\,
            I => \N__18716\
        );

    \I__4289\ : InMux
    port map (
            O => \N__18751\,
            I => \N__18709\
        );

    \I__4288\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18709\
        );

    \I__4287\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18709\
        );

    \I__4286\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18706\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__18745\,
            I => \N__18703\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__18742\,
            I => \N__18698\
        );

    \I__4283\ : Span4Mux_s3_v
    port map (
            O => \N__18739\,
            I => \N__18698\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__18736\,
            I => \N__18695\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__18731\,
            I => \N__18692\
        );

    \I__4280\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18689\
        );

    \I__4279\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18684\
        );

    \I__4278\ : InMux
    port map (
            O => \N__18728\,
            I => \N__18684\
        );

    \I__4277\ : Span4Mux_s3_h
    port map (
            O => \N__18725\,
            I => \N__18679\
        );

    \I__4276\ : Span4Mux_v
    port map (
            O => \N__18722\,
            I => \N__18679\
        );

    \I__4275\ : InMux
    port map (
            O => \N__18721\,
            I => \N__18672\
        );

    \I__4274\ : InMux
    port map (
            O => \N__18720\,
            I => \N__18672\
        );

    \I__4273\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18672\
        );

    \I__4272\ : Span4Mux_h
    port map (
            O => \N__18716\,
            I => \N__18667\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__18709\,
            I => \N__18667\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18658\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__18703\,
            I => \N__18658\
        );

    \I__4268\ : Span4Mux_v
    port map (
            O => \N__18698\,
            I => \N__18658\
        );

    \I__4267\ : Span4Mux_h
    port map (
            O => \N__18695\,
            I => \N__18658\
        );

    \I__4266\ : Odrv12
    port map (
            O => \N__18692\,
            I => \Lab_UT.un1_de_hex\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__18689\,
            I => \Lab_UT.un1_de_hex\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__18684\,
            I => \Lab_UT.un1_de_hex\
        );

    \I__4263\ : Odrv4
    port map (
            O => \N__18679\,
            I => \Lab_UT.un1_de_hex\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__18672\,
            I => \Lab_UT.un1_de_hex\
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__18667\,
            I => \Lab_UT.un1_de_hex\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__18658\,
            I => \Lab_UT.un1_de_hex\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__18643\,
            I => \N__18640\
        );

    \I__4258\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18637\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__18637\,
            I => \N__18634\
        );

    \I__4256\ : Span4Mux_s3_h
    port map (
            O => \N__18634\,
            I => \N__18631\
        );

    \I__4255\ : Odrv4
    port map (
            O => \N__18631\,
            I => \Lab_UT.scctrl.G_21_i_a7_0\
        );

    \I__4254\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18617\
        );

    \I__4253\ : CascadeMux
    port map (
            O => \N__18627\,
            I => \N__18613\
        );

    \I__4252\ : InMux
    port map (
            O => \N__18626\,
            I => \N__18608\
        );

    \I__4251\ : InMux
    port map (
            O => \N__18625\,
            I => \N__18605\
        );

    \I__4250\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18602\
        );

    \I__4249\ : InMux
    port map (
            O => \N__18623\,
            I => \N__18592\
        );

    \I__4248\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18592\
        );

    \I__4247\ : InMux
    port map (
            O => \N__18621\,
            I => \N__18592\
        );

    \I__4246\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18586\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__18617\,
            I => \N__18583\
        );

    \I__4244\ : InMux
    port map (
            O => \N__18616\,
            I => \N__18580\
        );

    \I__4243\ : InMux
    port map (
            O => \N__18613\,
            I => \N__18573\
        );

    \I__4242\ : InMux
    port map (
            O => \N__18612\,
            I => \N__18573\
        );

    \I__4241\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18573\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__18608\,
            I => \N__18566\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__18605\,
            I => \N__18566\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__18602\,
            I => \N__18563\
        );

    \I__4237\ : CascadeMux
    port map (
            O => \N__18601\,
            I => \N__18559\
        );

    \I__4236\ : CascadeMux
    port map (
            O => \N__18600\,
            I => \N__18556\
        );

    \I__4235\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18553\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__18592\,
            I => \N__18550\
        );

    \I__4233\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18547\
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__18590\,
            I => \N__18544\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__18589\,
            I => \N__18540\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__18586\,
            I => \N__18537\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__18583\,
            I => \N__18532\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__18580\,
            I => \N__18532\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__18573\,
            I => \N__18529\
        );

    \I__4226\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18524\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18524\
        );

    \I__4224\ : Span4Mux_v
    port map (
            O => \N__18566\,
            I => \N__18519\
        );

    \I__4223\ : Span4Mux_v
    port map (
            O => \N__18563\,
            I => \N__18519\
        );

    \I__4222\ : InMux
    port map (
            O => \N__18562\,
            I => \N__18512\
        );

    \I__4221\ : InMux
    port map (
            O => \N__18559\,
            I => \N__18512\
        );

    \I__4220\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18512\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__18553\,
            I => \N__18507\
        );

    \I__4218\ : Span4Mux_v
    port map (
            O => \N__18550\,
            I => \N__18507\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__18547\,
            I => \N__18504\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18497\
        );

    \I__4215\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18497\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18540\,
            I => \N__18497\
        );

    \I__4213\ : Span4Mux_h
    port map (
            O => \N__18537\,
            I => \N__18494\
        );

    \I__4212\ : Span4Mux_h
    port map (
            O => \N__18532\,
            I => \N__18491\
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__18529\,
            I => \Lab_UT.un4_de_hex\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__18524\,
            I => \Lab_UT.un4_de_hex\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__18519\,
            I => \Lab_UT.un4_de_hex\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__18512\,
            I => \Lab_UT.un4_de_hex\
        );

    \I__4207\ : Odrv4
    port map (
            O => \N__18507\,
            I => \Lab_UT.un4_de_hex\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__18504\,
            I => \Lab_UT.un4_de_hex\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__18497\,
            I => \Lab_UT.un4_de_hex\
        );

    \I__4204\ : Odrv4
    port map (
            O => \N__18494\,
            I => \Lab_UT.un4_de_hex\
        );

    \I__4203\ : Odrv4
    port map (
            O => \N__18491\,
            I => \Lab_UT.un4_de_hex\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__18472\,
            I => \Lab_UT.scctrl.g0_0_i_a8_0_1_cascade_\
        );

    \I__4201\ : InMux
    port map (
            O => \N__18469\,
            I => \N__18466\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__18466\,
            I => \N__18463\
        );

    \I__4199\ : Span4Mux_v
    port map (
            O => \N__18463\,
            I => \N__18460\
        );

    \I__4198\ : Span4Mux_h
    port map (
            O => \N__18460\,
            I => \N__18457\
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__18457\,
            I => \Lab_UT.scctrl.N_20\
        );

    \I__4196\ : CascadeMux
    port map (
            O => \N__18454\,
            I => \Lab_UT.scctrl.G_38_0_a3_0_4_cascade_\
        );

    \I__4195\ : InMux
    port map (
            O => \N__18451\,
            I => \N__18447\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__18450\,
            I => \N__18444\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__18447\,
            I => \N__18438\
        );

    \I__4192\ : InMux
    port map (
            O => \N__18444\,
            I => \N__18435\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__18443\,
            I => \N__18432\
        );

    \I__4190\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18429\
        );

    \I__4189\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18426\
        );

    \I__4188\ : Span4Mux_s1_h
    port map (
            O => \N__18438\,
            I => \N__18423\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__18435\,
            I => \N__18419\
        );

    \I__4186\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18416\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__18429\,
            I => \N__18413\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__18426\,
            I => \N__18410\
        );

    \I__4183\ : Span4Mux_v
    port map (
            O => \N__18423\,
            I => \N__18407\
        );

    \I__4182\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18404\
        );

    \I__4181\ : Span4Mux_s3_v
    port map (
            O => \N__18419\,
            I => \N__18399\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__18416\,
            I => \N__18399\
        );

    \I__4179\ : Span12Mux_s9_v
    port map (
            O => \N__18413\,
            I => \N__18396\
        );

    \I__4178\ : Span12Mux_s7_h
    port map (
            O => \N__18410\,
            I => \N__18393\
        );

    \I__4177\ : Odrv4
    port map (
            O => \N__18407\,
            I => \Lab_UT.scctrl.next_stateZ0Z_0\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__18404\,
            I => \Lab_UT.scctrl.next_stateZ0Z_0\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__18399\,
            I => \Lab_UT.scctrl.next_stateZ0Z_0\
        );

    \I__4174\ : Odrv12
    port map (
            O => \N__18396\,
            I => \Lab_UT.scctrl.next_stateZ0Z_0\
        );

    \I__4173\ : Odrv12
    port map (
            O => \N__18393\,
            I => \Lab_UT.scctrl.next_stateZ0Z_0\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__18382\,
            I => \Lab_UT.scctrl.G_38_0_1_cascade_\
        );

    \I__4171\ : InMux
    port map (
            O => \N__18379\,
            I => \N__18376\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__18376\,
            I => \Lab_UT.scctrl.N_7_0\
        );

    \I__4169\ : InMux
    port map (
            O => \N__18373\,
            I => \N__18370\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__18370\,
            I => \Lab_UT.scctrl.g0_0_i_0\
        );

    \I__4167\ : InMux
    port map (
            O => \N__18367\,
            I => \N__18364\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__18364\,
            I => \N__18361\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__18361\,
            I => \Lab_UT.scdp.a2b.g0_i_a9_1\
        );

    \I__4164\ : CascadeMux
    port map (
            O => \N__18358\,
            I => \Lab_UT.scdp.a2b.g0_iZ0Z_1_cascade_\
        );

    \I__4163\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18352\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__18352\,
            I => \N__18349\
        );

    \I__4161\ : Odrv12
    port map (
            O => \N__18349\,
            I => \Lab_UT.scdp.a2b.g0_iZ0Z_2\
        );

    \I__4160\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18343\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__18343\,
            I => \N__18340\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__18340\,
            I => \Lab_UT.scctrl.g1_i_a7_1\
        );

    \I__4157\ : CascadeMux
    port map (
            O => \N__18337\,
            I => \N__18333\
        );

    \I__4156\ : CascadeMux
    port map (
            O => \N__18336\,
            I => \N__18328\
        );

    \I__4155\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18322\
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__18332\,
            I => \N__18319\
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__18331\,
            I => \N__18316\
        );

    \I__4152\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18310\
        );

    \I__4151\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18310\
        );

    \I__4150\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18306\
        );

    \I__4149\ : InMux
    port map (
            O => \N__18325\,
            I => \N__18303\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__18322\,
            I => \N__18300\
        );

    \I__4147\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18293\
        );

    \I__4146\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18293\
        );

    \I__4145\ : InMux
    port map (
            O => \N__18315\,
            I => \N__18293\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__18310\,
            I => \N__18290\
        );

    \I__4143\ : InMux
    port map (
            O => \N__18309\,
            I => \N__18287\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__18306\,
            I => \N__18284\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__18303\,
            I => \N__18281\
        );

    \I__4140\ : Span4Mux_h
    port map (
            O => \N__18300\,
            I => \N__18276\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__18293\,
            I => \N__18276\
        );

    \I__4138\ : Span4Mux_h
    port map (
            O => \N__18290\,
            I => \N__18273\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__18287\,
            I => \N__18270\
        );

    \I__4136\ : Span4Mux_v
    port map (
            O => \N__18284\,
            I => \N__18263\
        );

    \I__4135\ : Span4Mux_h
    port map (
            O => \N__18281\,
            I => \N__18263\
        );

    \I__4134\ : Span4Mux_v
    port map (
            O => \N__18276\,
            I => \N__18263\
        );

    \I__4133\ : Span4Mux_v
    port map (
            O => \N__18273\,
            I => \N__18260\
        );

    \I__4132\ : Span4Mux_h
    port map (
            O => \N__18270\,
            I => \N__18257\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__18263\,
            I => \N__18254\
        );

    \I__4130\ : Odrv4
    port map (
            O => \N__18260\,
            I => \Lab_UT.scctrl.next_state_0_3\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__18257\,
            I => \Lab_UT.scctrl.next_state_0_3\
        );

    \I__4128\ : Odrv4
    port map (
            O => \N__18254\,
            I => \Lab_UT.scctrl.next_state_0_3\
        );

    \I__4127\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18243\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18240\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__18243\,
            I => \N__18237\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__18240\,
            I => \N__18231\
        );

    \I__4123\ : Span4Mux_v
    port map (
            O => \N__18237\,
            I => \N__18231\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18236\,
            I => \N__18228\
        );

    \I__4121\ : Odrv4
    port map (
            O => \N__18231\,
            I => \Lab_UT.scctrl.next_state_1_0_3\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__18228\,
            I => \Lab_UT.scctrl.next_state_1_0_3\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__18223\,
            I => \Lab_UT.scctrl.next_state_i_3_cascade_\
        );

    \I__4118\ : InMux
    port map (
            O => \N__18220\,
            I => \N__18217\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__18217\,
            I => \N__18213\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18216\,
            I => \N__18210\
        );

    \I__4115\ : Span4Mux_s3_v
    port map (
            O => \N__18213\,
            I => \N__18207\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__18210\,
            I => \N__18204\
        );

    \I__4113\ : Odrv4
    port map (
            O => \N__18207\,
            I => \Lab_UT.scctrl.next_state71\
        );

    \I__4112\ : Odrv4
    port map (
            O => \N__18204\,
            I => \Lab_UT.scctrl.next_state71\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18199\,
            I => \N__18195\
        );

    \I__4110\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18192\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__18195\,
            I => \N__18189\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__18192\,
            I => \N__18186\
        );

    \I__4107\ : Span4Mux_s3_v
    port map (
            O => \N__18189\,
            I => \N__18183\
        );

    \I__4106\ : Span4Mux_h
    port map (
            O => \N__18186\,
            I => \N__18180\
        );

    \I__4105\ : Odrv4
    port map (
            O => \N__18183\,
            I => \Lab_UT.scctrl.next_state72\
        );

    \I__4104\ : Odrv4
    port map (
            O => \N__18180\,
            I => \Lab_UT.scctrl.next_state72\
        );

    \I__4103\ : InMux
    port map (
            O => \N__18175\,
            I => \N__18172\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__18172\,
            I => \N__18169\
        );

    \I__4101\ : Odrv12
    port map (
            O => \N__18169\,
            I => \Lab_UT.scctrl.g4_1\
        );

    \I__4100\ : InMux
    port map (
            O => \N__18166\,
            I => \N__18157\
        );

    \I__4099\ : InMux
    port map (
            O => \N__18165\,
            I => \N__18157\
        );

    \I__4098\ : InMux
    port map (
            O => \N__18164\,
            I => \N__18157\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__18157\,
            I => \N__18152\
        );

    \I__4096\ : InMux
    port map (
            O => \N__18156\,
            I => \N__18147\
        );

    \I__4095\ : InMux
    port map (
            O => \N__18155\,
            I => \N__18147\
        );

    \I__4094\ : Span4Mux_v
    port map (
            O => \N__18152\,
            I => \N__18142\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__18147\,
            I => \N__18142\
        );

    \I__4092\ : Span4Mux_v
    port map (
            O => \N__18142\,
            I => \N__18137\
        );

    \I__4091\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18134\
        );

    \I__4090\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18131\
        );

    \I__4089\ : Span4Mux_h
    port map (
            O => \N__18137\,
            I => \N__18128\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__18134\,
            I => \N__18125\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18131\,
            I => \Lab_UT.sccEmsBitsSl\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__18128\,
            I => \Lab_UT.sccEmsBitsSl\
        );

    \I__4085\ : Odrv12
    port map (
            O => \N__18125\,
            I => \Lab_UT.sccEmsBitsSl\
        );

    \I__4084\ : InMux
    port map (
            O => \N__18118\,
            I => \N__18115\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__18115\,
            I => \N__18112\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__18112\,
            I => \Lab_UT.scctrl.g2\
        );

    \I__4081\ : InMux
    port map (
            O => \N__18109\,
            I => \N__18106\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__18106\,
            I => \N__18103\
        );

    \I__4079\ : Span4Mux_s3_v
    port map (
            O => \N__18103\,
            I => \N__18099\
        );

    \I__4078\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18096\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__18099\,
            I => \Lab_UT.scctrl.next_state_rst_3\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__18096\,
            I => \Lab_UT.scctrl.next_state_rst_3\
        );

    \I__4075\ : InMux
    port map (
            O => \N__18091\,
            I => \N__18088\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__18088\,
            I => \N__18035\
        );

    \I__4073\ : SRMux
    port map (
            O => \N__18087\,
            I => \N__17932\
        );

    \I__4072\ : SRMux
    port map (
            O => \N__18086\,
            I => \N__17932\
        );

    \I__4071\ : SRMux
    port map (
            O => \N__18085\,
            I => \N__17932\
        );

    \I__4070\ : SRMux
    port map (
            O => \N__18084\,
            I => \N__17932\
        );

    \I__4069\ : SRMux
    port map (
            O => \N__18083\,
            I => \N__17932\
        );

    \I__4068\ : SRMux
    port map (
            O => \N__18082\,
            I => \N__17932\
        );

    \I__4067\ : SRMux
    port map (
            O => \N__18081\,
            I => \N__17932\
        );

    \I__4066\ : SRMux
    port map (
            O => \N__18080\,
            I => \N__17932\
        );

    \I__4065\ : SRMux
    port map (
            O => \N__18079\,
            I => \N__17932\
        );

    \I__4064\ : SRMux
    port map (
            O => \N__18078\,
            I => \N__17932\
        );

    \I__4063\ : SRMux
    port map (
            O => \N__18077\,
            I => \N__17932\
        );

    \I__4062\ : SRMux
    port map (
            O => \N__18076\,
            I => \N__17932\
        );

    \I__4061\ : SRMux
    port map (
            O => \N__18075\,
            I => \N__17932\
        );

    \I__4060\ : SRMux
    port map (
            O => \N__18074\,
            I => \N__17932\
        );

    \I__4059\ : SRMux
    port map (
            O => \N__18073\,
            I => \N__17932\
        );

    \I__4058\ : SRMux
    port map (
            O => \N__18072\,
            I => \N__17932\
        );

    \I__4057\ : SRMux
    port map (
            O => \N__18071\,
            I => \N__17932\
        );

    \I__4056\ : SRMux
    port map (
            O => \N__18070\,
            I => \N__17932\
        );

    \I__4055\ : SRMux
    port map (
            O => \N__18069\,
            I => \N__17932\
        );

    \I__4054\ : SRMux
    port map (
            O => \N__18068\,
            I => \N__17932\
        );

    \I__4053\ : SRMux
    port map (
            O => \N__18067\,
            I => \N__17932\
        );

    \I__4052\ : SRMux
    port map (
            O => \N__18066\,
            I => \N__17932\
        );

    \I__4051\ : SRMux
    port map (
            O => \N__18065\,
            I => \N__17932\
        );

    \I__4050\ : SRMux
    port map (
            O => \N__18064\,
            I => \N__17932\
        );

    \I__4049\ : SRMux
    port map (
            O => \N__18063\,
            I => \N__17932\
        );

    \I__4048\ : SRMux
    port map (
            O => \N__18062\,
            I => \N__17932\
        );

    \I__4047\ : SRMux
    port map (
            O => \N__18061\,
            I => \N__17932\
        );

    \I__4046\ : SRMux
    port map (
            O => \N__18060\,
            I => \N__17932\
        );

    \I__4045\ : SRMux
    port map (
            O => \N__18059\,
            I => \N__17932\
        );

    \I__4044\ : SRMux
    port map (
            O => \N__18058\,
            I => \N__17932\
        );

    \I__4043\ : SRMux
    port map (
            O => \N__18057\,
            I => \N__17932\
        );

    \I__4042\ : SRMux
    port map (
            O => \N__18056\,
            I => \N__17932\
        );

    \I__4041\ : SRMux
    port map (
            O => \N__18055\,
            I => \N__17932\
        );

    \I__4040\ : SRMux
    port map (
            O => \N__18054\,
            I => \N__17932\
        );

    \I__4039\ : SRMux
    port map (
            O => \N__18053\,
            I => \N__17932\
        );

    \I__4038\ : SRMux
    port map (
            O => \N__18052\,
            I => \N__17932\
        );

    \I__4037\ : SRMux
    port map (
            O => \N__18051\,
            I => \N__17932\
        );

    \I__4036\ : SRMux
    port map (
            O => \N__18050\,
            I => \N__17932\
        );

    \I__4035\ : SRMux
    port map (
            O => \N__18049\,
            I => \N__17932\
        );

    \I__4034\ : SRMux
    port map (
            O => \N__18048\,
            I => \N__17932\
        );

    \I__4033\ : SRMux
    port map (
            O => \N__18047\,
            I => \N__17932\
        );

    \I__4032\ : SRMux
    port map (
            O => \N__18046\,
            I => \N__17932\
        );

    \I__4031\ : SRMux
    port map (
            O => \N__18045\,
            I => \N__17932\
        );

    \I__4030\ : SRMux
    port map (
            O => \N__18044\,
            I => \N__17932\
        );

    \I__4029\ : SRMux
    port map (
            O => \N__18043\,
            I => \N__17932\
        );

    \I__4028\ : SRMux
    port map (
            O => \N__18042\,
            I => \N__17932\
        );

    \I__4027\ : SRMux
    port map (
            O => \N__18041\,
            I => \N__17932\
        );

    \I__4026\ : SRMux
    port map (
            O => \N__18040\,
            I => \N__17932\
        );

    \I__4025\ : SRMux
    port map (
            O => \N__18039\,
            I => \N__17932\
        );

    \I__4024\ : SRMux
    port map (
            O => \N__18038\,
            I => \N__17932\
        );

    \I__4023\ : Glb2LocalMux
    port map (
            O => \N__18035\,
            I => \N__17932\
        );

    \I__4022\ : GlobalMux
    port map (
            O => \N__17932\,
            I => \N__17929\
        );

    \I__4021\ : gio2CtrlBuf
    port map (
            O => \N__17929\,
            I => \resetGen_rst_0_iso_g\
        );

    \I__4020\ : InMux
    port map (
            O => \N__17926\,
            I => \N__17922\
        );

    \I__4019\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17919\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__17922\,
            I => \N__17916\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__17919\,
            I => \N__17913\
        );

    \I__4016\ : Odrv12
    port map (
            O => \N__17916\,
            I => \Lab_UT.scctrl.next_state_rst_2\
        );

    \I__4015\ : Odrv4
    port map (
            O => \N__17913\,
            I => \Lab_UT.scctrl.next_state_rst_2\
        );

    \I__4014\ : InMux
    port map (
            O => \N__17908\,
            I => \N__17905\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__17905\,
            I => \Lab_UT.scctrl.N_223_2_reti\
        );

    \I__4012\ : InMux
    port map (
            O => \N__17902\,
            I => \N__17899\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__17899\,
            I => \N__17894\
        );

    \I__4010\ : InMux
    port map (
            O => \N__17898\,
            I => \N__17889\
        );

    \I__4009\ : InMux
    port map (
            O => \N__17897\,
            I => \N__17889\
        );

    \I__4008\ : Span4Mux_v
    port map (
            O => \N__17894\,
            I => \N__17883\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__17889\,
            I => \N__17883\
        );

    \I__4006\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17879\
        );

    \I__4005\ : Span4Mux_v
    port map (
            O => \N__17883\,
            I => \N__17876\
        );

    \I__4004\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17873\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__17879\,
            I => \N__17870\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__17876\,
            I => \Lab_UT.next_state_rst_2_0\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__17873\,
            I => \Lab_UT.next_state_rst_2_0\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__17870\,
            I => \Lab_UT.next_state_rst_2_0\
        );

    \I__3999\ : InMux
    port map (
            O => \N__17863\,
            I => \N__17860\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__17860\,
            I => \N__17857\
        );

    \I__3997\ : Span12Mux_s7_v
    port map (
            O => \N__17857\,
            I => \N__17854\
        );

    \I__3996\ : Odrv12
    port map (
            O => \N__17854\,
            I => \Lab_UT.scctrl.g0_i_3\
        );

    \I__3995\ : InMux
    port map (
            O => \N__17851\,
            I => \N__17848\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__17848\,
            I => \Lab_UT.scctrl.N_8\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__17845\,
            I => \Lab_UT.scctrl.g0_i_4_0_cascade_\
        );

    \I__3992\ : InMux
    port map (
            O => \N__17842\,
            I => \N__17833\
        );

    \I__3991\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17833\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__17840\,
            I => \N__17826\
        );

    \I__3989\ : InMux
    port map (
            O => \N__17839\,
            I => \N__17821\
        );

    \I__3988\ : InMux
    port map (
            O => \N__17838\,
            I => \N__17821\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__17833\,
            I => \N__17818\
        );

    \I__3986\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17811\
        );

    \I__3985\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17811\
        );

    \I__3984\ : InMux
    port map (
            O => \N__17830\,
            I => \N__17811\
        );

    \I__3983\ : InMux
    port map (
            O => \N__17829\,
            I => \N__17802\
        );

    \I__3982\ : InMux
    port map (
            O => \N__17826\,
            I => \N__17802\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__17821\,
            I => \N__17799\
        );

    \I__3980\ : Span4Mux_s3_v
    port map (
            O => \N__17818\,
            I => \N__17794\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__17811\,
            I => \N__17794\
        );

    \I__3978\ : InMux
    port map (
            O => \N__17810\,
            I => \N__17789\
        );

    \I__3977\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17789\
        );

    \I__3976\ : IoInMux
    port map (
            O => \N__17808\,
            I => \N__17786\
        );

    \I__3975\ : IoInMux
    port map (
            O => \N__17807\,
            I => \N__17783\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__17802\,
            I => \N__17780\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__17799\,
            I => \N__17773\
        );

    \I__3972\ : Span4Mux_v
    port map (
            O => \N__17794\,
            I => \N__17773\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__17789\,
            I => \N__17773\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__17786\,
            I => \N__17768\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__17783\,
            I => \N__17768\
        );

    \I__3968\ : Span4Mux_v
    port map (
            O => \N__17780\,
            I => \N__17765\
        );

    \I__3967\ : Span4Mux_h
    port map (
            O => \N__17773\,
            I => \N__17762\
        );

    \I__3966\ : Span4Mux_s0_h
    port map (
            O => \N__17768\,
            I => \N__17757\
        );

    \I__3965\ : Span4Mux_v
    port map (
            O => \N__17765\,
            I => \N__17757\
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__17762\,
            I => led_c_0
        );

    \I__3963\ : Odrv4
    port map (
            O => \N__17757\,
            I => led_c_0
        );

    \I__3962\ : InMux
    port map (
            O => \N__17752\,
            I => \N__17749\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__17749\,
            I => \N__17746\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__17746\,
            I => \Lab_UT.scctrl.N_8_1\
        );

    \I__3959\ : InMux
    port map (
            O => \N__17743\,
            I => \N__17740\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__17740\,
            I => \N__17737\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__17737\,
            I => \Lab_UT.scctrl.N_8_3\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__17734\,
            I => \Lab_UT.scctrl.g0_18_1_cascade_\
        );

    \I__3955\ : InMux
    port map (
            O => \N__17731\,
            I => \N__17727\
        );

    \I__3954\ : InMux
    port map (
            O => \N__17730\,
            I => \N__17724\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__17727\,
            I => \Lab_UT.scctrl.next_stateZ0Z_2\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__17724\,
            I => \Lab_UT.scctrl.next_stateZ0Z_2\
        );

    \I__3951\ : CascadeMux
    port map (
            O => \N__17719\,
            I => \Lab_UT.scctrl.next_stateZ0Z_2_cascade_\
        );

    \I__3950\ : InMux
    port map (
            O => \N__17716\,
            I => \N__17713\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__17713\,
            I => \Lab_UT.scctrl.N_6_2\
        );

    \I__3948\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17705\
        );

    \I__3947\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17700\
        );

    \I__3946\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17700\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__17705\,
            I => \Lab_UT.scctrl.g0_i_3_1\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__17700\,
            I => \Lab_UT.scctrl.g0_i_3_1\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__17695\,
            I => \N__17692\
        );

    \I__3942\ : InMux
    port map (
            O => \N__17692\,
            I => \N__17688\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__17691\,
            I => \N__17682\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__17688\,
            I => \N__17678\
        );

    \I__3939\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17675\
        );

    \I__3938\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17672\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__17685\,
            I => \N__17669\
        );

    \I__3936\ : InMux
    port map (
            O => \N__17682\,
            I => \N__17666\
        );

    \I__3935\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17663\
        );

    \I__3934\ : Span4Mux_s3_v
    port map (
            O => \N__17678\,
            I => \N__17660\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__17675\,
            I => \N__17655\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__17672\,
            I => \N__17655\
        );

    \I__3931\ : InMux
    port map (
            O => \N__17669\,
            I => \N__17652\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__17666\,
            I => \N__17645\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17663\,
            I => \N__17645\
        );

    \I__3928\ : Span4Mux_v
    port map (
            O => \N__17660\,
            I => \N__17645\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__17655\,
            I => next_state_1
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__17652\,
            I => next_state_1
        );

    \I__3925\ : Odrv4
    port map (
            O => \N__17645\,
            I => next_state_1
        );

    \I__3924\ : InMux
    port map (
            O => \N__17638\,
            I => \N__17635\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__17635\,
            I => \Lab_UT.scctrl.g0_i_m4_1_1\
        );

    \I__3922\ : InMux
    port map (
            O => \N__17632\,
            I => \N__17629\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__17629\,
            I => \Lab_UT.scctrl.N_9\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__17626\,
            I => \N__17620\
        );

    \I__3919\ : InMux
    port map (
            O => \N__17625\,
            I => \N__17617\
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__17624\,
            I => \N__17612\
        );

    \I__3917\ : InMux
    port map (
            O => \N__17623\,
            I => \N__17607\
        );

    \I__3916\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17604\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__17617\,
            I => \N__17601\
        );

    \I__3914\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17598\
        );

    \I__3913\ : CascadeMux
    port map (
            O => \N__17615\,
            I => \N__17595\
        );

    \I__3912\ : InMux
    port map (
            O => \N__17612\,
            I => \N__17590\
        );

    \I__3911\ : InMux
    port map (
            O => \N__17611\,
            I => \N__17590\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__17610\,
            I => \N__17587\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__17607\,
            I => \N__17584\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__17604\,
            I => \N__17577\
        );

    \I__3907\ : Span4Mux_h
    port map (
            O => \N__17601\,
            I => \N__17577\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__17598\,
            I => \N__17577\
        );

    \I__3905\ : InMux
    port map (
            O => \N__17595\,
            I => \N__17572\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__17590\,
            I => \N__17569\
        );

    \I__3903\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17566\
        );

    \I__3902\ : Span4Mux_v
    port map (
            O => \N__17584\,
            I => \N__17561\
        );

    \I__3901\ : Span4Mux_v
    port map (
            O => \N__17577\,
            I => \N__17561\
        );

    \I__3900\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17558\
        );

    \I__3899\ : InMux
    port map (
            O => \N__17575\,
            I => \N__17555\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__17572\,
            I => \N__17551\
        );

    \I__3897\ : Span4Mux_h
    port map (
            O => \N__17569\,
            I => \N__17540\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__17566\,
            I => \N__17540\
        );

    \I__3895\ : Span4Mux_h
    port map (
            O => \N__17561\,
            I => \N__17540\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__17558\,
            I => \N__17540\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__17555\,
            I => \N__17540\
        );

    \I__3892\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17537\
        );

    \I__3891\ : Span4Mux_h
    port map (
            O => \N__17551\,
            I => \N__17534\
        );

    \I__3890\ : Span4Mux_v
    port map (
            O => \N__17540\,
            I => \N__17531\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__17537\,
            I => rst_i_3_rep2
        );

    \I__3888\ : Odrv4
    port map (
            O => \N__17534\,
            I => rst_i_3_rep2
        );

    \I__3887\ : Odrv4
    port map (
            O => \N__17531\,
            I => rst_i_3_rep2
        );

    \I__3886\ : InMux
    port map (
            O => \N__17524\,
            I => \N__17521\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__17521\,
            I => \N__17517\
        );

    \I__3884\ : InMux
    port map (
            O => \N__17520\,
            I => \N__17514\
        );

    \I__3883\ : Odrv4
    port map (
            O => \N__17517\,
            I => \Lab_UT.state_ret_8_rep1_RNIJDTUE_1\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__17514\,
            I => \Lab_UT.state_ret_8_rep1_RNIJDTUE_1\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__17509\,
            I => \Lab_UT.scctrl.next_state_rst_0_5_0_cascade_\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__17506\,
            I => \N__17503\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17491\
        );

    \I__3878\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17486\
        );

    \I__3877\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17483\
        );

    \I__3876\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17477\
        );

    \I__3875\ : InMux
    port map (
            O => \N__17499\,
            I => \N__17477\
        );

    \I__3874\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17472\
        );

    \I__3873\ : InMux
    port map (
            O => \N__17497\,
            I => \N__17469\
        );

    \I__3872\ : InMux
    port map (
            O => \N__17496\,
            I => \N__17464\
        );

    \I__3871\ : InMux
    port map (
            O => \N__17495\,
            I => \N__17464\
        );

    \I__3870\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17461\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__17491\,
            I => \N__17458\
        );

    \I__3868\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17453\
        );

    \I__3867\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17453\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__17486\,
            I => \N__17450\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__17483\,
            I => \N__17447\
        );

    \I__3864\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17443\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__17477\,
            I => \N__17437\
        );

    \I__3862\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17432\
        );

    \I__3861\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17432\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__17472\,
            I => \N__17429\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__17469\,
            I => \N__17426\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__17464\,
            I => \N__17417\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__17461\,
            I => \N__17417\
        );

    \I__3856\ : Span4Mux_s3_h
    port map (
            O => \N__17458\,
            I => \N__17417\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__17453\,
            I => \N__17417\
        );

    \I__3854\ : Span4Mux_h
    port map (
            O => \N__17450\,
            I => \N__17412\
        );

    \I__3853\ : Span4Mux_v
    port map (
            O => \N__17447\,
            I => \N__17412\
        );

    \I__3852\ : InMux
    port map (
            O => \N__17446\,
            I => \N__17409\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__17443\,
            I => \N__17406\
        );

    \I__3850\ : InMux
    port map (
            O => \N__17442\,
            I => \N__17401\
        );

    \I__3849\ : InMux
    port map (
            O => \N__17441\,
            I => \N__17401\
        );

    \I__3848\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17398\
        );

    \I__3847\ : Span4Mux_h
    port map (
            O => \N__17437\,
            I => \N__17393\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__17432\,
            I => \N__17393\
        );

    \I__3845\ : Span12Mux_s4_v
    port map (
            O => \N__17429\,
            I => \N__17388\
        );

    \I__3844\ : Span12Mux_s11_v
    port map (
            O => \N__17426\,
            I => \N__17388\
        );

    \I__3843\ : Span4Mux_v
    port map (
            O => \N__17417\,
            I => \N__17383\
        );

    \I__3842\ : Span4Mux_v
    port map (
            O => \N__17412\,
            I => \N__17383\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__17409\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__3840\ : Odrv12
    port map (
            O => \N__17406\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__17401\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__17398\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__17393\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__3836\ : Odrv12
    port map (
            O => \N__17388\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__17383\,
            I => \Lab_UT.scctrl.stateZ0Z_3\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__17368\,
            I => \N__17364\
        );

    \I__3833\ : InMux
    port map (
            O => \N__17367\,
            I => \N__17360\
        );

    \I__3832\ : InMux
    port map (
            O => \N__17364\,
            I => \N__17356\
        );

    \I__3831\ : InMux
    port map (
            O => \N__17363\,
            I => \N__17353\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__17360\,
            I => \N__17350\
        );

    \I__3829\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17347\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__17356\,
            I => \N__17344\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__17353\,
            I => \N__17340\
        );

    \I__3826\ : Span4Mux_v
    port map (
            O => \N__17350\,
            I => \N__17337\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__17347\,
            I => \N__17333\
        );

    \I__3824\ : Span4Mux_h
    port map (
            O => \N__17344\,
            I => \N__17330\
        );

    \I__3823\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17327\
        );

    \I__3822\ : Span4Mux_h
    port map (
            O => \N__17340\,
            I => \N__17324\
        );

    \I__3821\ : Span4Mux_v
    port map (
            O => \N__17337\,
            I => \N__17321\
        );

    \I__3820\ : InMux
    port map (
            O => \N__17336\,
            I => \N__17318\
        );

    \I__3819\ : Span4Mux_h
    port map (
            O => \N__17333\,
            I => \N__17315\
        );

    \I__3818\ : Sp12to4
    port map (
            O => \N__17330\,
            I => \N__17310\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__17327\,
            I => \N__17310\
        );

    \I__3816\ : Odrv4
    port map (
            O => \N__17324\,
            I => rst_i_3_rep1
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__17321\,
            I => rst_i_3_rep1
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__17318\,
            I => rst_i_3_rep1
        );

    \I__3813\ : Odrv4
    port map (
            O => \N__17315\,
            I => rst_i_3_rep1
        );

    \I__3812\ : Odrv12
    port map (
            O => \N__17310\,
            I => rst_i_3_rep1
        );

    \I__3811\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17296\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__17296\,
            I => \Lab_UT.scctrl.g0_i_a8_1\
        );

    \I__3809\ : CascadeMux
    port map (
            O => \N__17293\,
            I => \N__17290\
        );

    \I__3808\ : InMux
    port map (
            O => \N__17290\,
            I => \N__17287\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__17287\,
            I => \Lab_UT.scctrl.g0_i_0_0\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17284\,
            I => \N__17281\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__17281\,
            I => \N__17278\
        );

    \I__3804\ : Odrv4
    port map (
            O => \N__17278\,
            I => \Lab_UT.scctrl.g0_7_3\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__17275\,
            I => \N__17272\
        );

    \I__3802\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17269\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__17269\,
            I => \Lab_UT.scctrl.g0_7_2\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__17266\,
            I => \Lab_UT.scctrl.g2_cascade_\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17263\,
            I => \N__17260\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__17260\,
            I => \Lab_UT.scctrl.g1_1\
        );

    \I__3797\ : InMux
    port map (
            O => \N__17257\,
            I => \N__17254\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__17254\,
            I => \N__17251\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__17251\,
            I => \Lab_UT.scctrl.g0_1_0\
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__17248\,
            I => \Lab_UT.scctrl.N_222i_cascade_\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17245\,
            I => \N__17242\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__17242\,
            I => \Lab_UT.scctrl.N_223_1_reti\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17239\,
            I => \N__17236\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__17236\,
            I => \N__17233\
        );

    \I__3789\ : Span4Mux_h
    port map (
            O => \N__17233\,
            I => \N__17230\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__17230\,
            I => \shifter_0_fast_RNI639J4_2\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__17227\,
            I => \Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433_cascade_\
        );

    \I__3786\ : InMux
    port map (
            O => \N__17224\,
            I => \N__17221\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17221\,
            I => \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17218\,
            I => \N__17212\
        );

    \I__3783\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17205\
        );

    \I__3782\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17205\
        );

    \I__3781\ : InMux
    port map (
            O => \N__17215\,
            I => \N__17205\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__17212\,
            I => \N__17202\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__17205\,
            I => \N__17199\
        );

    \I__3778\ : Span4Mux_v
    port map (
            O => \N__17202\,
            I => \N__17195\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__17199\,
            I => \N__17192\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17198\,
            I => \N__17189\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__17195\,
            I => \Lab_UT.de_bigD\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__17192\,
            I => \Lab_UT.de_bigD\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__17189\,
            I => \Lab_UT.de_bigD\
        );

    \I__3772\ : InMux
    port map (
            O => \N__17182\,
            I => \N__17179\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__17179\,
            I => \N__17175\
        );

    \I__3770\ : CascadeMux
    port map (
            O => \N__17178\,
            I => \N__17171\
        );

    \I__3769\ : Span4Mux_v
    port map (
            O => \N__17175\,
            I => \N__17167\
        );

    \I__3768\ : InMux
    port map (
            O => \N__17174\,
            I => \N__17160\
        );

    \I__3767\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17160\
        );

    \I__3766\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17160\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__17167\,
            I => \Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__17160\,
            I => \Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__17155\,
            I => \N__17151\
        );

    \I__3762\ : InMux
    port map (
            O => \N__17154\,
            I => \N__17145\
        );

    \I__3761\ : InMux
    port map (
            O => \N__17151\,
            I => \N__17136\
        );

    \I__3760\ : InMux
    port map (
            O => \N__17150\,
            I => \N__17136\
        );

    \I__3759\ : InMux
    port map (
            O => \N__17149\,
            I => \N__17136\
        );

    \I__3758\ : InMux
    port map (
            O => \N__17148\,
            I => \N__17136\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__17145\,
            I => \N__17132\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__17136\,
            I => \N__17129\
        );

    \I__3755\ : InMux
    port map (
            O => \N__17135\,
            I => \N__17126\
        );

    \I__3754\ : Odrv4
    port map (
            O => \N__17132\,
            I => \Lab_UT.de_bigL\
        );

    \I__3753\ : Odrv12
    port map (
            O => \N__17129\,
            I => \Lab_UT.de_bigL\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__17126\,
            I => \Lab_UT.de_bigL\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__17119\,
            I => \N__17116\
        );

    \I__3750\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17113\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__17113\,
            I => \N__17107\
        );

    \I__3748\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17100\
        );

    \I__3747\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17100\
        );

    \I__3746\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17100\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__17107\,
            I => \Lab_UT.scctrl.next_state_1_i_o2_0_d_1\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__17100\,
            I => \Lab_UT.scctrl.next_state_1_i_o2_0_d_1\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__17095\,
            I => \N__17092\
        );

    \I__3742\ : InMux
    port map (
            O => \N__17092\,
            I => \N__17086\
        );

    \I__3741\ : InMux
    port map (
            O => \N__17091\,
            I => \N__17086\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__17086\,
            I => \N__17083\
        );

    \I__3739\ : Span4Mux_v
    port map (
            O => \N__17083\,
            I => \N__17080\
        );

    \I__3738\ : Odrv4
    port map (
            O => \N__17080\,
            I => \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0Z_2\
        );

    \I__3737\ : InMux
    port map (
            O => \N__17077\,
            I => \N__17067\
        );

    \I__3736\ : InMux
    port map (
            O => \N__17076\,
            I => \N__17067\
        );

    \I__3735\ : InMux
    port map (
            O => \N__17075\,
            I => \N__17063\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17074\,
            I => \N__17060\
        );

    \I__3733\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17056\
        );

    \I__3732\ : InMux
    port map (
            O => \N__17072\,
            I => \N__17053\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__17067\,
            I => \N__17050\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17045\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17063\,
            I => \N__17042\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__17060\,
            I => \N__17039\
        );

    \I__3727\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17036\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__17056\,
            I => \N__17031\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__17053\,
            I => \N__17031\
        );

    \I__3724\ : Span4Mux_v
    port map (
            O => \N__17050\,
            I => \N__17028\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17023\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17048\,
            I => \N__17023\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__17045\,
            I => \N__17016\
        );

    \I__3720\ : Span4Mux_h
    port map (
            O => \N__17042\,
            I => \N__17011\
        );

    \I__3719\ : Span4Mux_h
    port map (
            O => \N__17039\,
            I => \N__17011\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__17036\,
            I => \N__17008\
        );

    \I__3717\ : Span4Mux_h
    port map (
            O => \N__17031\,
            I => \N__17005\
        );

    \I__3716\ : Span4Mux_s3_h
    port map (
            O => \N__17028\,
            I => \N__17002\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__17023\,
            I => \N__16999\
        );

    \I__3714\ : InMux
    port map (
            O => \N__17022\,
            I => \N__16994\
        );

    \I__3713\ : InMux
    port map (
            O => \N__17021\,
            I => \N__16994\
        );

    \I__3712\ : InMux
    port map (
            O => \N__17020\,
            I => \N__16989\
        );

    \I__3711\ : InMux
    port map (
            O => \N__17019\,
            I => \N__16989\
        );

    \I__3710\ : Odrv4
    port map (
            O => \N__17016\,
            I => bu_rx_data_6
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__17011\,
            I => bu_rx_data_6
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__17008\,
            I => bu_rx_data_6
        );

    \I__3707\ : Odrv4
    port map (
            O => \N__17005\,
            I => bu_rx_data_6
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__17002\,
            I => bu_rx_data_6
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__16999\,
            I => bu_rx_data_6
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__16994\,
            I => bu_rx_data_6
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__16989\,
            I => bu_rx_data_6
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__16972\,
            I => \N__16967\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__16971\,
            I => \N__16961\
        );

    \I__3700\ : InMux
    port map (
            O => \N__16970\,
            I => \N__16951\
        );

    \I__3699\ : InMux
    port map (
            O => \N__16967\,
            I => \N__16946\
        );

    \I__3698\ : InMux
    port map (
            O => \N__16966\,
            I => \N__16946\
        );

    \I__3697\ : InMux
    port map (
            O => \N__16965\,
            I => \N__16937\
        );

    \I__3696\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16934\
        );

    \I__3695\ : InMux
    port map (
            O => \N__16961\,
            I => \N__16931\
        );

    \I__3694\ : InMux
    port map (
            O => \N__16960\,
            I => \N__16928\
        );

    \I__3693\ : InMux
    port map (
            O => \N__16959\,
            I => \N__16921\
        );

    \I__3692\ : InMux
    port map (
            O => \N__16958\,
            I => \N__16921\
        );

    \I__3691\ : InMux
    port map (
            O => \N__16957\,
            I => \N__16921\
        );

    \I__3690\ : InMux
    port map (
            O => \N__16956\,
            I => \N__16918\
        );

    \I__3689\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16915\
        );

    \I__3688\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16912\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__16951\,
            I => \N__16909\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__16946\,
            I => \N__16906\
        );

    \I__3685\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16901\
        );

    \I__3684\ : InMux
    port map (
            O => \N__16944\,
            I => \N__16901\
        );

    \I__3683\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16896\
        );

    \I__3682\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16891\
        );

    \I__3681\ : InMux
    port map (
            O => \N__16941\,
            I => \N__16891\
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__16940\,
            I => \N__16887\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__16937\,
            I => \N__16883\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__16934\,
            I => \N__16880\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__16931\,
            I => \N__16874\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__16928\,
            I => \N__16867\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__16921\,
            I => \N__16867\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__16918\,
            I => \N__16867\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__16915\,
            I => \N__16864\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__16912\,
            I => \N__16855\
        );

    \I__3671\ : Span4Mux_v
    port map (
            O => \N__16909\,
            I => \N__16855\
        );

    \I__3670\ : Span4Mux_v
    port map (
            O => \N__16906\,
            I => \N__16855\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__16901\,
            I => \N__16855\
        );

    \I__3668\ : CascadeMux
    port map (
            O => \N__16900\,
            I => \N__16850\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__16899\,
            I => \N__16847\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__16896\,
            I => \N__16843\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__16891\,
            I => \N__16840\
        );

    \I__3664\ : InMux
    port map (
            O => \N__16890\,
            I => \N__16833\
        );

    \I__3663\ : InMux
    port map (
            O => \N__16887\,
            I => \N__16833\
        );

    \I__3662\ : InMux
    port map (
            O => \N__16886\,
            I => \N__16833\
        );

    \I__3661\ : Span4Mux_h
    port map (
            O => \N__16883\,
            I => \N__16828\
        );

    \I__3660\ : Span4Mux_h
    port map (
            O => \N__16880\,
            I => \N__16828\
        );

    \I__3659\ : InMux
    port map (
            O => \N__16879\,
            I => \N__16825\
        );

    \I__3658\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16820\
        );

    \I__3657\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16820\
        );

    \I__3656\ : Span4Mux_v
    port map (
            O => \N__16874\,
            I => \N__16815\
        );

    \I__3655\ : Span4Mux_v
    port map (
            O => \N__16867\,
            I => \N__16815\
        );

    \I__3654\ : Span4Mux_h
    port map (
            O => \N__16864\,
            I => \N__16810\
        );

    \I__3653\ : Span4Mux_h
    port map (
            O => \N__16855\,
            I => \N__16810\
        );

    \I__3652\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16801\
        );

    \I__3651\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16801\
        );

    \I__3650\ : InMux
    port map (
            O => \N__16850\,
            I => \N__16801\
        );

    \I__3649\ : InMux
    port map (
            O => \N__16847\,
            I => \N__16801\
        );

    \I__3648\ : InMux
    port map (
            O => \N__16846\,
            I => \N__16798\
        );

    \I__3647\ : Span4Mux_v
    port map (
            O => \N__16843\,
            I => \N__16791\
        );

    \I__3646\ : Span4Mux_v
    port map (
            O => \N__16840\,
            I => \N__16791\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__16833\,
            I => \N__16791\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__16828\,
            I => bu_rx_data_7
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__16825\,
            I => bu_rx_data_7
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__16820\,
            I => bu_rx_data_7
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__16815\,
            I => bu_rx_data_7
        );

    \I__3640\ : Odrv4
    port map (
            O => \N__16810\,
            I => bu_rx_data_7
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__16801\,
            I => bu_rx_data_7
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__16798\,
            I => bu_rx_data_7
        );

    \I__3637\ : Odrv4
    port map (
            O => \N__16791\,
            I => bu_rx_data_7
        );

    \I__3636\ : InMux
    port map (
            O => \N__16774\,
            I => \N__16771\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__16771\,
            I => \N__16768\
        );

    \I__3634\ : Span4Mux_v
    port map (
            O => \N__16768\,
            I => \N__16765\
        );

    \I__3633\ : Sp12to4
    port map (
            O => \N__16765\,
            I => \N__16762\
        );

    \I__3632\ : Odrv12
    port map (
            O => \N__16762\,
            I => \resetGen_escKey_4\
        );

    \I__3631\ : CEMux
    port map (
            O => \N__16759\,
            I => \N__16735\
        );

    \I__3630\ : CEMux
    port map (
            O => \N__16758\,
            I => \N__16735\
        );

    \I__3629\ : CEMux
    port map (
            O => \N__16757\,
            I => \N__16735\
        );

    \I__3628\ : CEMux
    port map (
            O => \N__16756\,
            I => \N__16735\
        );

    \I__3627\ : CEMux
    port map (
            O => \N__16755\,
            I => \N__16735\
        );

    \I__3626\ : CEMux
    port map (
            O => \N__16754\,
            I => \N__16735\
        );

    \I__3625\ : CEMux
    port map (
            O => \N__16753\,
            I => \N__16735\
        );

    \I__3624\ : CEMux
    port map (
            O => \N__16752\,
            I => \N__16735\
        );

    \I__3623\ : GlobalMux
    port map (
            O => \N__16735\,
            I => \N__16732\
        );

    \I__3622\ : gio2CtrlBuf
    port map (
            O => \N__16732\,
            I => \N_41_i_g\
        );

    \I__3621\ : InMux
    port map (
            O => \N__16729\,
            I => \N__16726\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__16726\,
            I => \N__16723\
        );

    \I__3619\ : Span4Mux_v
    port map (
            O => \N__16723\,
            I => \N__16720\
        );

    \I__3618\ : Span4Mux_s2_h
    port map (
            O => \N__16720\,
            I => \N__16717\
        );

    \I__3617\ : Span4Mux_h
    port map (
            O => \N__16717\,
            I => \N__16714\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__16714\,
            I => \Lab_UT.scctrl.g0_2_1\
        );

    \I__3615\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16708\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__16708\,
            I => \Lab_UT.scctrl.next_state_rst_0_3_N_6_0\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__16705\,
            I => \Lab_UT.scctrl.g1_0_0_cascade_\
        );

    \I__3612\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16699\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__16699\,
            I => \N__16696\
        );

    \I__3610\ : Odrv12
    port map (
            O => \N__16696\,
            I => \Lab_UT.scctrl.g0_1_3\
        );

    \I__3609\ : InMux
    port map (
            O => \N__16693\,
            I => \N__16690\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__16690\,
            I => \N__16687\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__16687\,
            I => \Lab_UT.scctrl.g0_1_0_0\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__16684\,
            I => \Lab_UT.scctrl.N_127_i_i_o6_0_1_cascade_\
        );

    \I__3605\ : InMux
    port map (
            O => \N__16681\,
            I => \N__16678\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__16678\,
            I => \Lab_UT.scctrl.N_127_i_i_a6_1\
        );

    \I__3603\ : InMux
    port map (
            O => \N__16675\,
            I => \N__16672\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__16672\,
            I => \Lab_UT.scctrl.N_190_0_0\
        );

    \I__3601\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16664\
        );

    \I__3600\ : InMux
    port map (
            O => \N__16668\,
            I => \N__16659\
        );

    \I__3599\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16659\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__16664\,
            I => \N__16656\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__16659\,
            I => \N__16653\
        );

    \I__3596\ : Span4Mux_h
    port map (
            O => \N__16656\,
            I => \N__16650\
        );

    \I__3595\ : Span4Mux_s3_h
    port map (
            O => \N__16653\,
            I => \N__16647\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__16650\,
            I => \Lab_UT.next_state_rst_0_5\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__16647\,
            I => \Lab_UT.next_state_rst_0_5\
        );

    \I__3592\ : InMux
    port map (
            O => \N__16642\,
            I => \N__16639\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__16639\,
            I => \Lab_UT.scdp.a2b.N_6_4\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__16636\,
            I => \N__16633\
        );

    \I__3589\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16630\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__16630\,
            I => \N__16627\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__16627\,
            I => \Lab_UT.state_ret_8_rep1_RNIHA8U3\
        );

    \I__3586\ : InMux
    port map (
            O => \N__16624\,
            I => \N__16618\
        );

    \I__3585\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16618\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__16618\,
            I => \Lab_UT.N_182\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16615\,
            I => \N__16612\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__16612\,
            I => \Lab_UT.scdp.a2b.g0_iZ0Z_9\
        );

    \I__3581\ : InMux
    port map (
            O => \N__16609\,
            I => \N__16606\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__16606\,
            I => \N__16600\
        );

    \I__3579\ : InMux
    port map (
            O => \N__16605\,
            I => \N__16593\
        );

    \I__3578\ : InMux
    port map (
            O => \N__16604\,
            I => \N__16593\
        );

    \I__3577\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16593\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__16600\,
            I => \Lab_UT.state_2_RNI3PVB9_2\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__16593\,
            I => \Lab_UT.state_2_RNI3PVB9_2\
        );

    \I__3574\ : InMux
    port map (
            O => \N__16588\,
            I => \N__16585\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__16585\,
            I => \Lab_UT.scctrl.N_182_0\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__16582\,
            I => \N__16578\
        );

    \I__3571\ : InMux
    port map (
            O => \N__16581\,
            I => \N__16575\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16578\,
            I => \N__16572\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__16575\,
            I => \N__16569\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__16572\,
            I => \N__16566\
        );

    \I__3567\ : Odrv12
    port map (
            O => \N__16569\,
            I => \Lab_UT.scctrl.N_166_0_1\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__16566\,
            I => \Lab_UT.scctrl.N_166_0_1\
        );

    \I__3565\ : InMux
    port map (
            O => \N__16561\,
            I => \N__16557\
        );

    \I__3564\ : InMux
    port map (
            O => \N__16560\,
            I => \N__16554\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__16557\,
            I => \N__16551\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__16554\,
            I => \N__16541\
        );

    \I__3561\ : Span4Mux_v
    port map (
            O => \N__16551\,
            I => \N__16541\
        );

    \I__3560\ : InMux
    port map (
            O => \N__16550\,
            I => \N__16538\
        );

    \I__3559\ : InMux
    port map (
            O => \N__16549\,
            I => \N__16535\
        );

    \I__3558\ : InMux
    port map (
            O => \N__16548\,
            I => \N__16532\
        );

    \I__3557\ : InMux
    port map (
            O => \N__16547\,
            I => \N__16527\
        );

    \I__3556\ : InMux
    port map (
            O => \N__16546\,
            I => \N__16527\
        );

    \I__3555\ : Span4Mux_h
    port map (
            O => \N__16541\,
            I => \N__16520\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__16538\,
            I => \N__16520\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__16535\,
            I => \N__16520\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__16532\,
            I => bu_rx_data_0_rep1
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__16527\,
            I => bu_rx_data_0_rep1
        );

    \I__3550\ : Odrv4
    port map (
            O => \N__16520\,
            I => bu_rx_data_0_rep1
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__16513\,
            I => \Lab_UT.scctrl.next_state_1_i_o2_0_d_1_cascade_\
        );

    \I__3548\ : InMux
    port map (
            O => \N__16510\,
            I => \N__16506\
        );

    \I__3547\ : InMux
    port map (
            O => \N__16509\,
            I => \N__16501\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__16506\,
            I => \N__16497\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__16505\,
            I => \N__16494\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__16504\,
            I => \N__16491\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__16501\,
            I => \N__16486\
        );

    \I__3542\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16483\
        );

    \I__3541\ : Span4Mux_h
    port map (
            O => \N__16497\,
            I => \N__16480\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16494\,
            I => \N__16477\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16491\,
            I => \N__16474\
        );

    \I__3538\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16471\
        );

    \I__3537\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16468\
        );

    \I__3536\ : Span4Mux_h
    port map (
            O => \N__16486\,
            I => \N__16463\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__16483\,
            I => \N__16463\
        );

    \I__3534\ : Odrv4
    port map (
            O => \N__16480\,
            I => \buart__rx_shifter_0_fast_2\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__16477\,
            I => \buart__rx_shifter_0_fast_2\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16474\,
            I => \buart__rx_shifter_0_fast_2\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__16471\,
            I => \buart__rx_shifter_0_fast_2\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__16468\,
            I => \buart__rx_shifter_0_fast_2\
        );

    \I__3529\ : Odrv4
    port map (
            O => \N__16463\,
            I => \buart__rx_shifter_0_fast_2\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__16450\,
            I => \Lab_UT.scctrl.next_state_rst_0_3_N_5L8Z0Z_1_cascade_\
        );

    \I__3527\ : InMux
    port map (
            O => \N__16447\,
            I => \N__16443\
        );

    \I__3526\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16440\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__16443\,
            I => \N__16437\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__16440\,
            I => \N__16434\
        );

    \I__3523\ : Span4Mux_v
    port map (
            O => \N__16437\,
            I => \N__16427\
        );

    \I__3522\ : Span4Mux_h
    port map (
            O => \N__16434\,
            I => \N__16427\
        );

    \I__3521\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16422\
        );

    \I__3520\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16422\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__16427\,
            I => \Lab_UT_dk_de_bigD_6\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__16422\,
            I => \Lab_UT_dk_de_bigD_6\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__16417\,
            I => \N__16414\
        );

    \I__3516\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16411\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__16411\,
            I => \Lab_UT.scctrl.g0_0_i_1_1\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__16408\,
            I => \N__16405\
        );

    \I__3513\ : InMux
    port map (
            O => \N__16405\,
            I => \N__16402\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__16402\,
            I => \N__16399\
        );

    \I__3511\ : Span4Mux_h
    port map (
            O => \N__16399\,
            I => \N__16396\
        );

    \I__3510\ : Odrv4
    port map (
            O => \N__16396\,
            I => \Lab_UT.scctrl.N_14\
        );

    \I__3509\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16390\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__16390\,
            I => \Lab_UT.scdp.a2b.g0_iZ0Z_4\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16387\,
            I => \N__16384\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__16384\,
            I => \Lab_UT.N_5\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__16381\,
            I => \Lab_UT.scdp.a2b.g0_iZ0Z_8_cascade_\
        );

    \I__3504\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16375\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__16375\,
            I => \Lab_UT.scdp.a2b.g0_3_a3_6\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__16372\,
            I => \N__16368\
        );

    \I__3501\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16364\
        );

    \I__3500\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16359\
        );

    \I__3499\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16359\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__16364\,
            I => \N__16355\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__16359\,
            I => \N__16349\
        );

    \I__3496\ : InMux
    port map (
            O => \N__16358\,
            I => \N__16346\
        );

    \I__3495\ : Span4Mux_v
    port map (
            O => \N__16355\,
            I => \N__16343\
        );

    \I__3494\ : InMux
    port map (
            O => \N__16354\,
            I => \N__16338\
        );

    \I__3493\ : InMux
    port map (
            O => \N__16353\,
            I => \N__16333\
        );

    \I__3492\ : InMux
    port map (
            O => \N__16352\,
            I => \N__16333\
        );

    \I__3491\ : Span4Mux_v
    port map (
            O => \N__16349\,
            I => \N__16330\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__16346\,
            I => \N__16327\
        );

    \I__3489\ : Span4Mux_s2_h
    port map (
            O => \N__16343\,
            I => \N__16324\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16342\,
            I => \N__16319\
        );

    \I__3487\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16319\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__16338\,
            I => \Lab_UT.de_cr_2\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__16333\,
            I => \Lab_UT.de_cr_2\
        );

    \I__3484\ : Odrv4
    port map (
            O => \N__16330\,
            I => \Lab_UT.de_cr_2\
        );

    \I__3483\ : Odrv4
    port map (
            O => \N__16327\,
            I => \Lab_UT.de_cr_2\
        );

    \I__3482\ : Odrv4
    port map (
            O => \N__16324\,
            I => \Lab_UT.de_cr_2\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__16319\,
            I => \Lab_UT.de_cr_2\
        );

    \I__3480\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16301\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16298\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__16304\,
            I => \N__16294\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__16301\,
            I => \N__16286\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__16298\,
            I => \N__16286\
        );

    \I__3475\ : InMux
    port map (
            O => \N__16297\,
            I => \N__16283\
        );

    \I__3474\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16280\
        );

    \I__3473\ : CascadeMux
    port map (
            O => \N__16293\,
            I => \N__16277\
        );

    \I__3472\ : CascadeMux
    port map (
            O => \N__16292\,
            I => \N__16274\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__16291\,
            I => \N__16271\
        );

    \I__3470\ : Span4Mux_v
    port map (
            O => \N__16286\,
            I => \N__16267\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__16283\,
            I => \N__16264\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__16280\,
            I => \N__16261\
        );

    \I__3467\ : InMux
    port map (
            O => \N__16277\,
            I => \N__16256\
        );

    \I__3466\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16256\
        );

    \I__3465\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16251\
        );

    \I__3464\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16251\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__16267\,
            I => \Lab_UT.de_cr_6_0\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__16264\,
            I => \Lab_UT.de_cr_6_0\
        );

    \I__3461\ : Odrv12
    port map (
            O => \N__16261\,
            I => \Lab_UT.de_cr_6_0\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__16256\,
            I => \Lab_UT.de_cr_6_0\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__16251\,
            I => \Lab_UT.de_cr_6_0\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__16240\,
            I => \Lab_UT.g0_i_a5_1_3_cascade_\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16237\,
            I => \N__16234\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__16234\,
            I => \Lab_UT.scdp.a2b.N_9_1\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__16231\,
            I => \N__16227\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__16230\,
            I => \N__16224\
        );

    \I__3453\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16221\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16218\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__16221\,
            I => \Lab_UT.scdp.a2b.g1_1_0_1\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__16218\,
            I => \Lab_UT.scdp.a2b.g1_1_0_1\
        );

    \I__3449\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16210\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__16210\,
            I => \Lab_UT.scctrl.g0_1_3_1\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16207\,
            I => \N__16204\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__16204\,
            I => \N__16201\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__16201\,
            I => \N__16198\
        );

    \I__3444\ : Span4Mux_s3_h
    port map (
            O => \N__16198\,
            I => \N__16195\
        );

    \I__3443\ : Odrv4
    port map (
            O => \N__16195\,
            I => \Lab_UT_dk_de_cr_12_1\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__16192\,
            I => \N__16189\
        );

    \I__3441\ : InMux
    port map (
            O => \N__16189\,
            I => \N__16186\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__16186\,
            I => \N__16181\
        );

    \I__3439\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16176\
        );

    \I__3438\ : InMux
    port map (
            O => \N__16184\,
            I => \N__16176\
        );

    \I__3437\ : Odrv12
    port map (
            O => \N__16181\,
            I => \ufifo.emptyB_0\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__16176\,
            I => \ufifo.emptyB_0\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__16171\,
            I => \N__16159\
        );

    \I__3434\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16156\
        );

    \I__3433\ : InMux
    port map (
            O => \N__16169\,
            I => \N__16150\
        );

    \I__3432\ : InMux
    port map (
            O => \N__16168\,
            I => \N__16150\
        );

    \I__3431\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16147\
        );

    \I__3430\ : InMux
    port map (
            O => \N__16166\,
            I => \N__16143\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16137\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16164\,
            I => \N__16137\
        );

    \I__3427\ : InMux
    port map (
            O => \N__16163\,
            I => \N__16133\
        );

    \I__3426\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16128\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16128\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__16156\,
            I => \N__16125\
        );

    \I__3423\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16122\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__16150\,
            I => \N__16119\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__16147\,
            I => \N__16116\
        );

    \I__3420\ : InMux
    port map (
            O => \N__16146\,
            I => \N__16113\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__16143\,
            I => \N__16110\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16142\,
            I => \N__16107\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__16137\,
            I => \N__16104\
        );

    \I__3416\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16101\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__16133\,
            I => \N__16096\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__16128\,
            I => \N__16096\
        );

    \I__3413\ : Span4Mux_h
    port map (
            O => \N__16125\,
            I => \N__16089\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__16122\,
            I => \N__16089\
        );

    \I__3411\ : Span4Mux_h
    port map (
            O => \N__16119\,
            I => \N__16089\
        );

    \I__3410\ : Span4Mux_h
    port map (
            O => \N__16116\,
            I => \N__16076\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__16113\,
            I => \N__16076\
        );

    \I__3408\ : Span4Mux_h
    port map (
            O => \N__16110\,
            I => \N__16076\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__16107\,
            I => \N__16076\
        );

    \I__3406\ : Span4Mux_h
    port map (
            O => \N__16104\,
            I => \N__16076\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__16101\,
            I => \N__16076\
        );

    \I__3404\ : Odrv4
    port map (
            O => \N__16096\,
            I => bu_rx_data_0
        );

    \I__3403\ : Odrv4
    port map (
            O => \N__16089\,
            I => bu_rx_data_0
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__16076\,
            I => bu_rx_data_0
        );

    \I__3401\ : InMux
    port map (
            O => \N__16069\,
            I => \N__16066\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__16066\,
            I => \N__16063\
        );

    \I__3399\ : Odrv12
    port map (
            O => \N__16063\,
            I => \ufifo.tx_fsm.N_60_0\
        );

    \I__3398\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16057\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__16057\,
            I => \N__16054\
        );

    \I__3396\ : Span4Mux_h
    port map (
            O => \N__16054\,
            I => \N__16051\
        );

    \I__3395\ : Odrv4
    port map (
            O => \N__16051\,
            I => \Lab_UT.scctrl.N_127_i_i_a6_0_0\
        );

    \I__3394\ : InMux
    port map (
            O => \N__16048\,
            I => \N__16045\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__16045\,
            I => \Lab_UT.scctrl.N_11\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16042\,
            I => \N__16039\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__16039\,
            I => \Lab_UT.scctrl.G_21_i_a7_1_1\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__16036\,
            I => \N__16033\
        );

    \I__3389\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16030\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__16030\,
            I => \N__16027\
        );

    \I__3387\ : Odrv12
    port map (
            O => \N__16027\,
            I => \Lab_UT.m61_i_a2_2\
        );

    \I__3386\ : InMux
    port map (
            O => \N__16024\,
            I => \N__16021\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__16021\,
            I => \Lab_UT.scctrl.g0_0_i_0_0\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__16018\,
            I => \Lab_UT.N_5_cascade_\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16015\,
            I => \N__16012\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__16012\,
            I => \Lab_UT.g0_i_5\
        );

    \I__3381\ : InMux
    port map (
            O => \N__16009\,
            I => \N__16006\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__16006\,
            I => \Lab_UT.scctrl.g0_14_mb_sn\
        );

    \I__3379\ : InMux
    port map (
            O => \N__16003\,
            I => \N__16000\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__16000\,
            I => \G_23_0_0\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__15997\,
            I => \N__15994\
        );

    \I__3376\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15991\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__15991\,
            I => \N__15988\
        );

    \I__3374\ : Odrv4
    port map (
            O => \N__15988\,
            I => \Lab_UT.scctrl.N_12_1\
        );

    \I__3373\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15981\
        );

    \I__3372\ : InMux
    port map (
            O => \N__15984\,
            I => \N__15978\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__15981\,
            I => \Lab_UT.scctrl.N_5_0\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__15978\,
            I => \Lab_UT.scctrl.N_5_0\
        );

    \I__3369\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15970\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__15970\,
            I => \N__15967\
        );

    \I__3367\ : Odrv4
    port map (
            O => \N__15967\,
            I => \Lab_UT.scctrl.g0_0_i_a8_3_1_0\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__15964\,
            I => \Lab_UT.scctrl.g0_0_i_a8_2_1_0_cascade_\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__15961\,
            I => \Lab_UT.scctrl.g0_0_i_3_0_cascade_\
        );

    \I__3364\ : InMux
    port map (
            O => \N__15958\,
            I => \N__15955\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__15955\,
            I => \Lab_UT.scctrl.N_13\
        );

    \I__3362\ : InMux
    port map (
            O => \N__15952\,
            I => \N__15949\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__15949\,
            I => \Lab_UT.scctrl.g0_i_1\
        );

    \I__3360\ : InMux
    port map (
            O => \N__15946\,
            I => \N__15936\
        );

    \I__3359\ : InMux
    port map (
            O => \N__15945\,
            I => \N__15936\
        );

    \I__3358\ : InMux
    port map (
            O => \N__15944\,
            I => \N__15936\
        );

    \I__3357\ : InMux
    port map (
            O => \N__15943\,
            I => \N__15933\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__15936\,
            I => \Lab_UT.scctrl.g0_0_i_2\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__15933\,
            I => \Lab_UT.scctrl.g0_0_i_2\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__15928\,
            I => \N__15925\
        );

    \I__3353\ : InMux
    port map (
            O => \N__15925\,
            I => \N__15915\
        );

    \I__3352\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15915\
        );

    \I__3351\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15915\
        );

    \I__3350\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15911\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__15915\,
            I => \N__15908\
        );

    \I__3348\ : InMux
    port map (
            O => \N__15914\,
            I => \N__15905\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__15911\,
            I => \Lab_UT.scctrl.g0_16_mb_sn\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__15908\,
            I => \Lab_UT.scctrl.g0_16_mb_sn\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__15905\,
            I => \Lab_UT.scctrl.g0_16_mb_sn\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__15898\,
            I => \N__15892\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__15897\,
            I => \N__15888\
        );

    \I__3342\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15885\
        );

    \I__3341\ : InMux
    port map (
            O => \N__15895\,
            I => \N__15878\
        );

    \I__3340\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15878\
        );

    \I__3339\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15878\
        );

    \I__3338\ : InMux
    port map (
            O => \N__15888\,
            I => \N__15875\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__15885\,
            I => \N__15868\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__15878\,
            I => \N__15868\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__15875\,
            I => \N__15868\
        );

    \I__3334\ : Span4Mux_v
    port map (
            O => \N__15868\,
            I => \N__15865\
        );

    \I__3333\ : Span4Mux_s3_h
    port map (
            O => \N__15865\,
            I => \N__15862\
        );

    \I__3332\ : Odrv4
    port map (
            O => \N__15862\,
            I => \Lab_UT.scctrl.g0_16_mb_rn_0\
        );

    \I__3331\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15853\
        );

    \I__3330\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15848\
        );

    \I__3329\ : InMux
    port map (
            O => \N__15857\,
            I => \N__15848\
        );

    \I__3328\ : InMux
    port map (
            O => \N__15856\,
            I => \N__15845\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__15853\,
            I => \Lab_UT.scctrl.g0_0_i_3_0\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__15848\,
            I => \Lab_UT.scctrl.g0_0_i_3_0\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__15845\,
            I => \Lab_UT.scctrl.g0_0_i_3_0\
        );

    \I__3324\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15835\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__15835\,
            I => \N__15831\
        );

    \I__3322\ : InMux
    port map (
            O => \N__15834\,
            I => \N__15828\
        );

    \I__3321\ : Span4Mux_h
    port map (
            O => \N__15831\,
            I => \N__15825\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__15828\,
            I => \Lab_UT.scdp.key0_5\
        );

    \I__3319\ : Odrv4
    port map (
            O => \N__15825\,
            I => \Lab_UT.scdp.key0_5\
        );

    \I__3318\ : InMux
    port map (
            O => \N__15820\,
            I => \N__15813\
        );

    \I__3317\ : InMux
    port map (
            O => \N__15819\,
            I => \N__15813\
        );

    \I__3316\ : InMux
    port map (
            O => \N__15818\,
            I => \N__15810\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__15813\,
            I => \N__15806\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__15810\,
            I => \N__15803\
        );

    \I__3313\ : InMux
    port map (
            O => \N__15809\,
            I => \N__15800\
        );

    \I__3312\ : Span4Mux_h
    port map (
            O => \N__15806\,
            I => \N__15793\
        );

    \I__3311\ : Span4Mux_h
    port map (
            O => \N__15803\,
            I => \N__15793\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__15800\,
            I => \N__15793\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__15793\,
            I => \Lab_UT.scdp.a2b.N_53\
        );

    \I__3308\ : CascadeMux
    port map (
            O => \N__15790\,
            I => \N__15786\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__15789\,
            I => \N__15783\
        );

    \I__3306\ : InMux
    port map (
            O => \N__15786\,
            I => \N__15777\
        );

    \I__3305\ : InMux
    port map (
            O => \N__15783\,
            I => \N__15777\
        );

    \I__3304\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15773\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__15777\,
            I => \N__15768\
        );

    \I__3302\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15765\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__15773\,
            I => \N__15762\
        );

    \I__3300\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15759\
        );

    \I__3299\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15755\
        );

    \I__3298\ : Span4Mux_h
    port map (
            O => \N__15768\,
            I => \N__15747\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__15765\,
            I => \N__15747\
        );

    \I__3296\ : Span4Mux_v
    port map (
            O => \N__15762\,
            I => \N__15742\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__15759\,
            I => \N__15742\
        );

    \I__3294\ : InMux
    port map (
            O => \N__15758\,
            I => \N__15739\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__15755\,
            I => \N__15736\
        );

    \I__3292\ : InMux
    port map (
            O => \N__15754\,
            I => \N__15733\
        );

    \I__3291\ : InMux
    port map (
            O => \N__15753\,
            I => \N__15728\
        );

    \I__3290\ : InMux
    port map (
            O => \N__15752\,
            I => \N__15728\
        );

    \I__3289\ : Span4Mux_v
    port map (
            O => \N__15747\,
            I => \N__15723\
        );

    \I__3288\ : Span4Mux_h
    port map (
            O => \N__15742\,
            I => \N__15723\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__15739\,
            I => \N__15720\
        );

    \I__3286\ : Span4Mux_v
    port map (
            O => \N__15736\,
            I => \N__15717\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__15733\,
            I => bu_rx_data_1
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__15728\,
            I => bu_rx_data_1
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__15723\,
            I => bu_rx_data_1
        );

    \I__3282\ : Odrv12
    port map (
            O => \N__15720\,
            I => bu_rx_data_1
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__15717\,
            I => bu_rx_data_1
        );

    \I__3280\ : InMux
    port map (
            O => \N__15706\,
            I => \N__15697\
        );

    \I__3279\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15697\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__15704\,
            I => \N__15691\
        );

    \I__3277\ : CascadeMux
    port map (
            O => \N__15703\,
            I => \N__15688\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__15702\,
            I => \N__15683\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__15697\,
            I => \N__15677\
        );

    \I__3274\ : InMux
    port map (
            O => \N__15696\,
            I => \N__15674\
        );

    \I__3273\ : InMux
    port map (
            O => \N__15695\,
            I => \N__15671\
        );

    \I__3272\ : InMux
    port map (
            O => \N__15694\,
            I => \N__15666\
        );

    \I__3271\ : InMux
    port map (
            O => \N__15691\,
            I => \N__15666\
        );

    \I__3270\ : InMux
    port map (
            O => \N__15688\,
            I => \N__15662\
        );

    \I__3269\ : InMux
    port map (
            O => \N__15687\,
            I => \N__15659\
        );

    \I__3268\ : InMux
    port map (
            O => \N__15686\,
            I => \N__15656\
        );

    \I__3267\ : InMux
    port map (
            O => \N__15683\,
            I => \N__15653\
        );

    \I__3266\ : InMux
    port map (
            O => \N__15682\,
            I => \N__15647\
        );

    \I__3265\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15642\
        );

    \I__3264\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15642\
        );

    \I__3263\ : Span4Mux_v
    port map (
            O => \N__15677\,
            I => \N__15639\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__15674\,
            I => \N__15636\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__15671\,
            I => \N__15633\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__15666\,
            I => \N__15630\
        );

    \I__3259\ : InMux
    port map (
            O => \N__15665\,
            I => \N__15627\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__15662\,
            I => \N__15624\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__15659\,
            I => \N__15621\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__15656\,
            I => \N__15618\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__15653\,
            I => \N__15615\
        );

    \I__3254\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15612\
        );

    \I__3253\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15607\
        );

    \I__3252\ : InMux
    port map (
            O => \N__15650\,
            I => \N__15607\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__15647\,
            I => \N__15602\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__15642\,
            I => \N__15602\
        );

    \I__3249\ : Span4Mux_v
    port map (
            O => \N__15639\,
            I => \N__15593\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__15636\,
            I => \N__15593\
        );

    \I__3247\ : Span4Mux_v
    port map (
            O => \N__15633\,
            I => \N__15593\
        );

    \I__3246\ : Span4Mux_v
    port map (
            O => \N__15630\,
            I => \N__15593\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__15627\,
            I => \N__15588\
        );

    \I__3244\ : Span4Mux_h
    port map (
            O => \N__15624\,
            I => \N__15588\
        );

    \I__3243\ : Span4Mux_v
    port map (
            O => \N__15621\,
            I => \N__15581\
        );

    \I__3242\ : Span4Mux_v
    port map (
            O => \N__15618\,
            I => \N__15581\
        );

    \I__3241\ : Span4Mux_s2_h
    port map (
            O => \N__15615\,
            I => \N__15581\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__15612\,
            I => bu_rx_data_2
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__15607\,
            I => bu_rx_data_2
        );

    \I__3238\ : Odrv12
    port map (
            O => \N__15602\,
            I => bu_rx_data_2
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__15593\,
            I => bu_rx_data_2
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__15588\,
            I => bu_rx_data_2
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__15581\,
            I => bu_rx_data_2
        );

    \I__3234\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15562\
        );

    \I__3233\ : InMux
    port map (
            O => \N__15567\,
            I => \N__15562\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__15562\,
            I => \N__15553\
        );

    \I__3231\ : InMux
    port map (
            O => \N__15561\,
            I => \N__15550\
        );

    \I__3230\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15541\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15541\
        );

    \I__3228\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15541\
        );

    \I__3227\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15541\
        );

    \I__3226\ : InMux
    port map (
            O => \N__15556\,
            I => \N__15538\
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__15553\,
            I => \Lab_UT.scdp.binValD_2\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15550\,
            I => \Lab_UT.scdp.binValD_2\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__15541\,
            I => \Lab_UT.scdp.binValD_2\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__15538\,
            I => \Lab_UT.scdp.binValD_2\
        );

    \I__3221\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15525\
        );

    \I__3220\ : InMux
    port map (
            O => \N__15528\,
            I => \N__15522\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__15525\,
            I => \N__15519\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__15522\,
            I => \N__15514\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__15519\,
            I => \N__15514\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__15514\,
            I => \Lab_UT.scdp.key0_6\
        );

    \I__3215\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15506\
        );

    \I__3214\ : InMux
    port map (
            O => \N__15510\,
            I => \N__15503\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__15509\,
            I => \N__15500\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__15506\,
            I => \N__15494\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__15503\,
            I => \N__15491\
        );

    \I__3210\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15482\
        );

    \I__3209\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15482\
        );

    \I__3208\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15482\
        );

    \I__3207\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15479\
        );

    \I__3206\ : Span4Mux_v
    port map (
            O => \N__15494\,
            I => \N__15474\
        );

    \I__3205\ : Span4Mux_v
    port map (
            O => \N__15491\,
            I => \N__15474\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15469\
        );

    \I__3203\ : InMux
    port map (
            O => \N__15489\,
            I => \N__15469\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__15482\,
            I => \N__15464\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__15479\,
            I => \N__15464\
        );

    \I__3200\ : Span4Mux_s3_h
    port map (
            O => \N__15474\,
            I => \N__15461\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__15469\,
            I => \Lab_UT.scdp.binValD_0\
        );

    \I__3198\ : Odrv12
    port map (
            O => \N__15464\,
            I => \Lab_UT.scdp.binValD_0\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__15461\,
            I => \Lab_UT.scdp.binValD_0\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15454\,
            I => \N__15451\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__15451\,
            I => \N__15448\
        );

    \I__3194\ : Span4Mux_v
    port map (
            O => \N__15448\,
            I => \N__15444\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15447\,
            I => \N__15441\
        );

    \I__3192\ : Span4Mux_s2_v
    port map (
            O => \N__15444\,
            I => \N__15438\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__15441\,
            I => \Lab_UT.scdp.key0_4\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__15438\,
            I => \Lab_UT.scdp.key0_4\
        );

    \I__3189\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15426\
        );

    \I__3188\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15417\
        );

    \I__3187\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15417\
        );

    \I__3186\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15417\
        );

    \I__3185\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15417\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__15426\,
            I => \Lab_UT.state_ret_RNIUV0941_0\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__15417\,
            I => \Lab_UT.state_ret_RNIUV0941_0\
        );

    \I__3182\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15408\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__15411\,
            I => \N__15405\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__15408\,
            I => \N__15402\
        );

    \I__3179\ : InMux
    port map (
            O => \N__15405\,
            I => \N__15399\
        );

    \I__3178\ : Span4Mux_h
    port map (
            O => \N__15402\,
            I => \N__15396\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__15399\,
            I => \Lab_UT.scdp.key0_7\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__15396\,
            I => \Lab_UT.scdp.key0_7\
        );

    \I__3175\ : CascadeMux
    port map (
            O => \N__15391\,
            I => \N__15387\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__15390\,
            I => \N__15380\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15369\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15386\,
            I => \N__15369\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15385\,
            I => \N__15369\
        );

    \I__3170\ : InMux
    port map (
            O => \N__15384\,
            I => \N__15369\
        );

    \I__3169\ : InMux
    port map (
            O => \N__15383\,
            I => \N__15369\
        );

    \I__3168\ : InMux
    port map (
            O => \N__15380\,
            I => \N__15366\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__15369\,
            I => \N__15361\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__15366\,
            I => \N__15358\
        );

    \I__3165\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15353\
        );

    \I__3164\ : InMux
    port map (
            O => \N__15364\,
            I => \N__15353\
        );

    \I__3163\ : Span4Mux_s2_v
    port map (
            O => \N__15361\,
            I => \N__15350\
        );

    \I__3162\ : Odrv12
    port map (
            O => \N__15358\,
            I => \Lab_UT.scdp.binValD_1\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__15353\,
            I => \Lab_UT.scdp.binValD_1\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__15350\,
            I => \Lab_UT.scdp.binValD_1\
        );

    \I__3159\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15340\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__15340\,
            I => \N__15336\
        );

    \I__3157\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15333\
        );

    \I__3156\ : Span4Mux_h
    port map (
            O => \N__15336\,
            I => \N__15330\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__15333\,
            I => \Lab_UT.scdp.key0_1\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__15330\,
            I => \Lab_UT.scdp.key0_1\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15318\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15313\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15323\,
            I => \N__15306\
        );

    \I__3150\ : InMux
    port map (
            O => \N__15322\,
            I => \N__15306\
        );

    \I__3149\ : InMux
    port map (
            O => \N__15321\,
            I => \N__15306\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__15318\,
            I => \N__15303\
        );

    \I__3147\ : InMux
    port map (
            O => \N__15317\,
            I => \N__15298\
        );

    \I__3146\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15298\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__15313\,
            I => \N__15291\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__15306\,
            I => \N__15291\
        );

    \I__3143\ : Span4Mux_s2_v
    port map (
            O => \N__15303\,
            I => \N__15291\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__15298\,
            I => \Lab_UT.scdp.binValD_3\
        );

    \I__3141\ : Odrv4
    port map (
            O => \N__15291\,
            I => \Lab_UT.scdp.binValD_3\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__15286\,
            I => \N__15283\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15283\,
            I => \N__15269\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__15282\,
            I => \N__15266\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__15281\,
            I => \N__15262\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__15280\,
            I => \N__15259\
        );

    \I__3135\ : CascadeMux
    port map (
            O => \N__15279\,
            I => \N__15256\
        );

    \I__3134\ : CascadeMux
    port map (
            O => \N__15278\,
            I => \N__15253\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__15277\,
            I => \N__15244\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__15276\,
            I => \N__15241\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__15275\,
            I => \N__15237\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__15274\,
            I => \N__15234\
        );

    \I__3129\ : CascadeMux
    port map (
            O => \N__15273\,
            I => \N__15225\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__15272\,
            I => \N__15220\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__15269\,
            I => \N__15217\
        );

    \I__3126\ : InMux
    port map (
            O => \N__15266\,
            I => \N__15214\
        );

    \I__3125\ : InMux
    port map (
            O => \N__15265\,
            I => \N__15203\
        );

    \I__3124\ : InMux
    port map (
            O => \N__15262\,
            I => \N__15203\
        );

    \I__3123\ : InMux
    port map (
            O => \N__15259\,
            I => \N__15203\
        );

    \I__3122\ : InMux
    port map (
            O => \N__15256\,
            I => \N__15203\
        );

    \I__3121\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15203\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__15252\,
            I => \N__15200\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__15251\,
            I => \N__15197\
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__15250\,
            I => \N__15194\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__15249\,
            I => \N__15191\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__15248\,
            I => \N__15188\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__15247\,
            I => \N__15185\
        );

    \I__3114\ : InMux
    port map (
            O => \N__15244\,
            I => \N__15175\
        );

    \I__3113\ : InMux
    port map (
            O => \N__15241\,
            I => \N__15175\
        );

    \I__3112\ : InMux
    port map (
            O => \N__15240\,
            I => \N__15175\
        );

    \I__3111\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15158\
        );

    \I__3110\ : InMux
    port map (
            O => \N__15234\,
            I => \N__15158\
        );

    \I__3109\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15158\
        );

    \I__3108\ : InMux
    port map (
            O => \N__15232\,
            I => \N__15158\
        );

    \I__3107\ : InMux
    port map (
            O => \N__15231\,
            I => \N__15158\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15158\
        );

    \I__3105\ : InMux
    port map (
            O => \N__15229\,
            I => \N__15158\
        );

    \I__3104\ : InMux
    port map (
            O => \N__15228\,
            I => \N__15158\
        );

    \I__3103\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15151\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15224\,
            I => \N__15151\
        );

    \I__3101\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15151\
        );

    \I__3100\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15148\
        );

    \I__3099\ : Span4Mux_v
    port map (
            O => \N__15217\,
            I => \N__15143\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__15214\,
            I => \N__15143\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__15203\,
            I => \N__15140\
        );

    \I__3096\ : InMux
    port map (
            O => \N__15200\,
            I => \N__15135\
        );

    \I__3095\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15135\
        );

    \I__3094\ : InMux
    port map (
            O => \N__15194\,
            I => \N__15132\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15129\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15118\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15185\,
            I => \N__15118\
        );

    \I__3090\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15118\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15118\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15118\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__15175\,
            I => \N__15115\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__15158\,
            I => \N__15112\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__15151\,
            I => \N__15109\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__15148\,
            I => \N__15104\
        );

    \I__3083\ : Span4Mux_h
    port map (
            O => \N__15143\,
            I => \N__15104\
        );

    \I__3082\ : Span4Mux_h
    port map (
            O => \N__15140\,
            I => \N__15101\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__15135\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__15132\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__15129\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__15118\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__15115\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__3076\ : Odrv12
    port map (
            O => \N__15112\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__3075\ : Odrv12
    port map (
            O => \N__15109\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__3074\ : Odrv4
    port map (
            O => \N__15104\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__15101\,
            I => \Lab_UT.scdp.binVal_ValidD\
        );

    \I__3072\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15078\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15072\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__15078\,
            I => \N__15069\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15066\
        );

    \I__3068\ : InMux
    port map (
            O => \N__15076\,
            I => \N__15061\
        );

    \I__3067\ : InMux
    port map (
            O => \N__15075\,
            I => \N__15061\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__15072\,
            I => \Lab_UT.state_0_RNIKFK051_0_1\
        );

    \I__3065\ : Odrv4
    port map (
            O => \N__15069\,
            I => \Lab_UT.state_0_RNIKFK051_0_1\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__15066\,
            I => \Lab_UT.state_0_RNIKFK051_0_1\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__15061\,
            I => \Lab_UT.state_0_RNIKFK051_0_1\
        );

    \I__3062\ : InMux
    port map (
            O => \N__15052\,
            I => \N__15049\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__15049\,
            I => \N__15045\
        );

    \I__3060\ : InMux
    port map (
            O => \N__15048\,
            I => \N__15042\
        );

    \I__3059\ : Span4Mux_h
    port map (
            O => \N__15045\,
            I => \N__15039\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__15042\,
            I => \Lab_UT.scdp.key0_3\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__15039\,
            I => \Lab_UT.scdp.key0_3\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15034\,
            I => \N__15031\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__15031\,
            I => \N__15027\
        );

    \I__3054\ : InMux
    port map (
            O => \N__15030\,
            I => \N__15024\
        );

    \I__3053\ : Span4Mux_v
    port map (
            O => \N__15027\,
            I => \N__15021\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__15024\,
            I => \N__15018\
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__15021\,
            I => \Lab_UT.scctrl.next_state74\
        );

    \I__3050\ : Odrv4
    port map (
            O => \N__15018\,
            I => \Lab_UT.scctrl.next_state74\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__15013\,
            I => \N__15010\
        );

    \I__3048\ : InMux
    port map (
            O => \N__15010\,
            I => \N__15007\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__15007\,
            I => \N__15004\
        );

    \I__3046\ : Odrv12
    port map (
            O => \N__15004\,
            I => \Lab_UT.scctrl.N_7_1\
        );

    \I__3045\ : InMux
    port map (
            O => \N__15001\,
            I => \N__14998\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__14998\,
            I => \Lab_UT.scctrl.N_223_2\
        );

    \I__3043\ : InMux
    port map (
            O => \N__14995\,
            I => \N__14992\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__14992\,
            I => \Lab_UT.scctrl.next_state73\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__14989\,
            I => \Lab_UT.scctrl.next_state73_cascade_\
        );

    \I__3040\ : InMux
    port map (
            O => \N__14986\,
            I => \N__14973\
        );

    \I__3039\ : InMux
    port map (
            O => \N__14985\,
            I => \N__14973\
        );

    \I__3038\ : InMux
    port map (
            O => \N__14984\,
            I => \N__14973\
        );

    \I__3037\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14970\
        );

    \I__3036\ : InMux
    port map (
            O => \N__14982\,
            I => \N__14967\
        );

    \I__3035\ : InMux
    port map (
            O => \N__14981\,
            I => \N__14964\
        );

    \I__3034\ : InMux
    port map (
            O => \N__14980\,
            I => \N__14961\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__14973\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__14970\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__14967\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__14964\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__14961\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__14950\,
            I => \Lab_UT.state_ret_3_RNII68F41_0_cascade_\
        );

    \I__3027\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14944\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__14944\,
            I => \N__14940\
        );

    \I__3025\ : InMux
    port map (
            O => \N__14943\,
            I => \N__14937\
        );

    \I__3024\ : Span4Mux_h
    port map (
            O => \N__14940\,
            I => \N__14934\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__14937\,
            I => \Lab_UT.scdp.key2_0\
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__14934\,
            I => \Lab_UT.scdp.key2_0\
        );

    \I__3021\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14925\
        );

    \I__3020\ : InMux
    port map (
            O => \N__14928\,
            I => \N__14922\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__14925\,
            I => \N__14919\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__14922\,
            I => \N__14914\
        );

    \I__3017\ : Span4Mux_h
    port map (
            O => \N__14919\,
            I => \N__14914\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__14914\,
            I => \Lab_UT.scdp.key2_1\
        );

    \I__3015\ : InMux
    port map (
            O => \N__14911\,
            I => \N__14905\
        );

    \I__3014\ : InMux
    port map (
            O => \N__14910\,
            I => \N__14898\
        );

    \I__3013\ : InMux
    port map (
            O => \N__14909\,
            I => \N__14898\
        );

    \I__3012\ : InMux
    port map (
            O => \N__14908\,
            I => \N__14898\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__14905\,
            I => \Lab_UT.state_ret_3_RNII68F41_0\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__14898\,
            I => \Lab_UT.state_ret_3_RNII68F41_0\
        );

    \I__3009\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14890\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__14890\,
            I => \N__14887\
        );

    \I__3007\ : Span4Mux_v
    port map (
            O => \N__14887\,
            I => \N__14883\
        );

    \I__3006\ : InMux
    port map (
            O => \N__14886\,
            I => \N__14880\
        );

    \I__3005\ : Span4Mux_h
    port map (
            O => \N__14883\,
            I => \N__14877\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__14880\,
            I => \Lab_UT.scdp.key2_2\
        );

    \I__3003\ : Odrv4
    port map (
            O => \N__14877\,
            I => \Lab_UT.scdp.key2_2\
        );

    \I__3002\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14869\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__14869\,
            I => \N__14863\
        );

    \I__3000\ : InMux
    port map (
            O => \N__14868\,
            I => \N__14856\
        );

    \I__2999\ : InMux
    port map (
            O => \N__14867\,
            I => \N__14856\
        );

    \I__2998\ : InMux
    port map (
            O => \N__14866\,
            I => \N__14856\
        );

    \I__2997\ : Span4Mux_v
    port map (
            O => \N__14863\,
            I => \N__14849\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__14856\,
            I => \N__14849\
        );

    \I__2995\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14846\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__14854\,
            I => \N__14841\
        );

    \I__2993\ : Span4Mux_h
    port map (
            O => \N__14849\,
            I => \N__14838\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__14846\,
            I => \N__14835\
        );

    \I__2991\ : InMux
    port map (
            O => \N__14845\,
            I => \N__14830\
        );

    \I__2990\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14830\
        );

    \I__2989\ : InMux
    port map (
            O => \N__14841\,
            I => \N__14827\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__14838\,
            I => bu_rx_data_i_3_1
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__14835\,
            I => bu_rx_data_i_3_1
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__14830\,
            I => bu_rx_data_i_3_1
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__14827\,
            I => bu_rx_data_i_3_1
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__14818\,
            I => \N__14815\
        );

    \I__2983\ : InMux
    port map (
            O => \N__14815\,
            I => \N__14809\
        );

    \I__2982\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14809\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__14809\,
            I => \Lab_UT.scctrl.g0_i_2_0\
        );

    \I__2980\ : InMux
    port map (
            O => \N__14806\,
            I => \N__14802\
        );

    \I__2979\ : InMux
    port map (
            O => \N__14805\,
            I => \N__14799\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__14802\,
            I => \Lab_UT.scctrl.next_state_rst_0_3_N_6_1\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__14799\,
            I => \Lab_UT.scctrl.next_state_rst_0_3_N_6_1\
        );

    \I__2976\ : CEMux
    port map (
            O => \N__14794\,
            I => \N__14788\
        );

    \I__2975\ : CEMux
    port map (
            O => \N__14793\,
            I => \N__14785\
        );

    \I__2974\ : CEMux
    port map (
            O => \N__14792\,
            I => \N__14782\
        );

    \I__2973\ : CEMux
    port map (
            O => \N__14791\,
            I => \N__14779\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__14788\,
            I => \N__14776\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__14785\,
            I => \N__14773\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__14782\,
            I => \N__14770\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__14779\,
            I => \N__14767\
        );

    \I__2968\ : Span4Mux_v
    port map (
            O => \N__14776\,
            I => \N__14762\
        );

    \I__2967\ : Span4Mux_h
    port map (
            O => \N__14773\,
            I => \N__14762\
        );

    \I__2966\ : Span4Mux_v
    port map (
            O => \N__14770\,
            I => \N__14757\
        );

    \I__2965\ : Span4Mux_v
    port map (
            O => \N__14767\,
            I => \N__14757\
        );

    \I__2964\ : Odrv4
    port map (
            O => \N__14762\,
            I => \Lab_UT.g0_3_0\
        );

    \I__2963\ : Odrv4
    port map (
            O => \N__14757\,
            I => \Lab_UT.g0_3_0\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__14752\,
            I => \N__14749\
        );

    \I__2961\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14746\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__14746\,
            I => \Lab_UT.scctrl.g0_i_a8_3_0\
        );

    \I__2959\ : InMux
    port map (
            O => \N__14743\,
            I => \N__14740\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__14740\,
            I => \Lab_UT.scctrl.N_6_3\
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__14737\,
            I => \Lab_UT.scctrl.g0_i_1_1_cascade_\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__14734\,
            I => \Lab_UT.scctrl.next_state_1_0_1_3_cascade_\
        );

    \I__2955\ : InMux
    port map (
            O => \N__14731\,
            I => \N__14728\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__14728\,
            I => \N__14724\
        );

    \I__2953\ : InMux
    port map (
            O => \N__14727\,
            I => \N__14721\
        );

    \I__2952\ : Odrv4
    port map (
            O => \N__14724\,
            I => \Lab_UT.scctrl.next_state75\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__14721\,
            I => \Lab_UT.scctrl.next_state75\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__14716\,
            I => \Lab_UT.scctrl.next_state_rst_1_3_1_cascade_\
        );

    \I__2949\ : InMux
    port map (
            O => \N__14713\,
            I => \N__14710\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__14710\,
            I => \N__14707\
        );

    \I__2947\ : Odrv4
    port map (
            O => \N__14707\,
            I => \Lab_UT.next_state_rst_1_3\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__14704\,
            I => \Lab_UT.next_state_rst_1_3_cascade_\
        );

    \I__2945\ : InMux
    port map (
            O => \N__14701\,
            I => \N__14697\
        );

    \I__2944\ : InMux
    port map (
            O => \N__14700\,
            I => \N__14694\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__14697\,
            I => \N__14691\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__14694\,
            I => \N__14688\
        );

    \I__2941\ : Span4Mux_h
    port map (
            O => \N__14691\,
            I => \N__14685\
        );

    \I__2940\ : Odrv12
    port map (
            O => \N__14688\,
            I => \Lab_UT.scctrl.N_166_0\
        );

    \I__2939\ : Odrv4
    port map (
            O => \N__14685\,
            I => \Lab_UT.scctrl.N_166_0\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__14680\,
            I => \Lab_UT.scctrl.next_state_rst_1_cascade_\
        );

    \I__2937\ : CascadeMux
    port map (
            O => \N__14677\,
            I => \N__14673\
        );

    \I__2936\ : InMux
    port map (
            O => \N__14676\,
            I => \N__14669\
        );

    \I__2935\ : InMux
    port map (
            O => \N__14673\,
            I => \N__14666\
        );

    \I__2934\ : IoInMux
    port map (
            O => \N__14672\,
            I => \N__14663\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__14669\,
            I => \N__14660\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__14666\,
            I => \N__14657\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__14663\,
            I => \N__14654\
        );

    \I__2930\ : Span4Mux_v
    port map (
            O => \N__14660\,
            I => \N__14651\
        );

    \I__2929\ : Span4Mux_h
    port map (
            O => \N__14657\,
            I => \N__14648\
        );

    \I__2928\ : Odrv12
    port map (
            O => \N__14654\,
            I => led_c_2
        );

    \I__2927\ : Odrv4
    port map (
            O => \N__14651\,
            I => led_c_2
        );

    \I__2926\ : Odrv4
    port map (
            O => \N__14648\,
            I => led_c_2
        );

    \I__2925\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14638\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__14638\,
            I => \N__14635\
        );

    \I__2923\ : Span4Mux_v
    port map (
            O => \N__14635\,
            I => \N__14632\
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__14632\,
            I => \Lab_UT.scctrl.g0_17_N_4LZ0Z5\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__14629\,
            I => \Lab_UT.scctrl.next_state_rst_0_3_N_6_1_cascade_\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__14626\,
            I => \Lab_UT.scctrl.g0_i_2_0_cascade_\
        );

    \I__2919\ : InMux
    port map (
            O => \N__14623\,
            I => \N__14617\
        );

    \I__2918\ : InMux
    port map (
            O => \N__14622\,
            I => \N__14617\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__14617\,
            I => \Lab_UT.scctrl.next_state_rst_0\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__14614\,
            I => \Lab_UT.scctrl.g0_1_1_cascade_\
        );

    \I__2915\ : InMux
    port map (
            O => \N__14611\,
            I => \N__14608\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__14608\,
            I => \Lab_UT.scctrl.g0_2_0\
        );

    \I__2913\ : InMux
    port map (
            O => \N__14605\,
            I => \N__14602\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__14602\,
            I => \N__14599\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__14599\,
            I => \Lab_UT.scctrl.N_12_0\
        );

    \I__2910\ : InMux
    port map (
            O => \N__14596\,
            I => \N__14593\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__14593\,
            I => \Lab_UT.scctrl.g0_i_1_0\
        );

    \I__2908\ : CascadeMux
    port map (
            O => \N__14590\,
            I => \Lab_UT.scctrl.g0_i_3_0_cascade_\
        );

    \I__2907\ : InMux
    port map (
            O => \N__14587\,
            I => \N__14584\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__14584\,
            I => \N__14581\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__14581\,
            I => \Lab_UT.scctrl.un6_sccDecrypt_0\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__14578\,
            I => \Lab_UT.scctrl.g1_1_0_cascade_\
        );

    \I__2903\ : InMux
    port map (
            O => \N__14575\,
            I => \N__14572\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__14572\,
            I => \Lab_UT.scctrl.g2_0\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__14569\,
            I => \Lab_UT.scctrl.g0_1_2_cascade_\
        );

    \I__2900\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14563\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__14563\,
            I => \Lab_UT.scctrl.g0_8_0\
        );

    \I__2898\ : InMux
    port map (
            O => \N__14560\,
            I => \N__14557\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__14557\,
            I => \Lab_UT.scdp.a2b.g1_1_o2_0Z0Z_0\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__14554\,
            I => \Lab_UT.scdp.a2b.N_6_1_cascade_\
        );

    \I__2895\ : InMux
    port map (
            O => \N__14551\,
            I => \N__14548\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__14548\,
            I => \Lab_UT.scdp.a2b.g0_3_a3_0Z0Z_3\
        );

    \I__2893\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14542\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__14542\,
            I => \N__14539\
        );

    \I__2891\ : Span4Mux_h
    port map (
            O => \N__14539\,
            I => \N__14533\
        );

    \I__2890\ : InMux
    port map (
            O => \N__14538\,
            I => \N__14526\
        );

    \I__2889\ : InMux
    port map (
            O => \N__14537\,
            I => \N__14526\
        );

    \I__2888\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14526\
        );

    \I__2887\ : Odrv4
    port map (
            O => \N__14533\,
            I => \Lab_UT.N_190\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__14526\,
            I => \Lab_UT.N_190\
        );

    \I__2885\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14518\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__14518\,
            I => \N__14515\
        );

    \I__2883\ : Span4Mux_h
    port map (
            O => \N__14515\,
            I => \N__14512\
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__14512\,
            I => \Lab_UT.scctrl.N_6_3_0\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__14509\,
            I => \N_127_i_i_1_cascade_\
        );

    \I__2880\ : InMux
    port map (
            O => \N__14506\,
            I => \N__14503\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__14503\,
            I => \N__14500\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__14500\,
            I => \Lab_UT.scctrl.N_11_0\
        );

    \I__2877\ : InMux
    port map (
            O => \N__14497\,
            I => \N__14494\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__14494\,
            I => \Lab_UT.N_166_0_0\
        );

    \I__2875\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14488\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__14488\,
            I => \Lab_UT.scctrl.N_127_i_i_3\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__14485\,
            I => \Lab_UT.g1_i_a4_0_2_cascade_\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__14482\,
            I => \N__14479\
        );

    \I__2871\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14476\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__14476\,
            I => \N__14470\
        );

    \I__2869\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14467\
        );

    \I__2868\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14464\
        );

    \I__2867\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14461\
        );

    \I__2866\ : Span4Mux_v
    port map (
            O => \N__14470\,
            I => \N__14452\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__14467\,
            I => \N__14452\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__14464\,
            I => \N__14452\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__14461\,
            I => \N__14452\
        );

    \I__2862\ : Odrv4
    port map (
            O => \N__14452\,
            I => \Lab_UT.next_state_3\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__14449\,
            I => \Lab_UT.g0_3_a3_0_4_cascade_\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__14446\,
            I => \Lab_UT.scctrl.g0_0_i_2_cascade_\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__14443\,
            I => \N__14439\
        );

    \I__2858\ : InMux
    port map (
            O => \N__14442\,
            I => \N__14434\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14439\,
            I => \N__14434\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__14434\,
            I => \N__14430\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14433\,
            I => \N__14427\
        );

    \I__2854\ : Span4Mux_h
    port map (
            O => \N__14430\,
            I => \N__14424\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__14427\,
            I => \N__14421\
        );

    \I__2852\ : Span4Mux_v
    port map (
            O => \N__14424\,
            I => \N__14418\
        );

    \I__2851\ : Span4Mux_v
    port map (
            O => \N__14421\,
            I => \N__14415\
        );

    \I__2850\ : Odrv4
    port map (
            O => \N__14418\,
            I => \Lab_UT.scctrl.state_i_3_fast_0\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__14415\,
            I => \Lab_UT.scctrl.state_i_3_fast_0\
        );

    \I__2848\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14407\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__14407\,
            I => \Lab_UT.scctrl.g0_i_1_1_0\
        );

    \I__2846\ : InMux
    port map (
            O => \N__14404\,
            I => \N__14401\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__14401\,
            I => \N__14398\
        );

    \I__2844\ : Span4Mux_h
    port map (
            O => \N__14398\,
            I => \N__14395\
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__14395\,
            I => \Lab_UT.scdp.a2b.N_6_0\
        );

    \I__2842\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14389\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__14389\,
            I => \N__14386\
        );

    \I__2840\ : Span4Mux_v
    port map (
            O => \N__14386\,
            I => \N__14383\
        );

    \I__2839\ : Span4Mux_s3_h
    port map (
            O => \N__14383\,
            I => \N__14380\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__14380\,
            I => \Lab_UT.scctrl.g0_14_mb_rn_0\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__14377\,
            I => \Lab_UT.scctrl.g0_0_i_1_cascade_\
        );

    \I__2836\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14371\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__14371\,
            I => \Lab_UT.scctrl.N_7_2\
        );

    \I__2834\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14365\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__14365\,
            I => \N__14362\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__14362\,
            I => \Lab_UT.scctrl.state_i_3_fast_2\
        );

    \I__2831\ : InMux
    port map (
            O => \N__14359\,
            I => \N__14356\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__14356\,
            I => \N__14353\
        );

    \I__2829\ : Span4Mux_h
    port map (
            O => \N__14353\,
            I => \N__14350\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__14350\,
            I => \Lab_UT.scctrl.next_state_1_0_a5_0_0_3\
        );

    \I__2827\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14343\
        );

    \I__2826\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14340\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14343\,
            I => \Lab_UT.scctrl.g0_i_4\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__14340\,
            I => \Lab_UT.scctrl.g0_i_4\
        );

    \I__2823\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14332\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__14332\,
            I => \N__14328\
        );

    \I__2821\ : InMux
    port map (
            O => \N__14331\,
            I => \N__14325\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__14328\,
            I => \Lab_UT.scctrl.N_10\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__14325\,
            I => \Lab_UT.scctrl.N_10\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__14320\,
            I => \Lab_UT.scctrl.G_23_0_a9_4_2_cascade_\
        );

    \I__2817\ : InMux
    port map (
            O => \N__14317\,
            I => \N__14314\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__14314\,
            I => \Lab_UT.scctrl.G_23_0_3\
        );

    \I__2815\ : InMux
    port map (
            O => \N__14311\,
            I => \N__14305\
        );

    \I__2814\ : InMux
    port map (
            O => \N__14310\,
            I => \N__14305\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__14305\,
            I => \Lab_UT.scctrl.G_23_0_a9_3_1\
        );

    \I__2812\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14296\
        );

    \I__2811\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14296\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__14296\,
            I => \Lab_UT.scctrl.G_23_0_4\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__14293\,
            I => \Lab_UT.scctrl.G_23_0_3_cascade_\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14290\,
            I => \N__14286\
        );

    \I__2807\ : InMux
    port map (
            O => \N__14289\,
            I => \N__14283\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__14286\,
            I => \Lab_UT.scctrl.N_3ctr\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__14283\,
            I => \Lab_UT.scctrl.N_3ctr\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__14278\,
            I => \N__14275\
        );

    \I__2803\ : InMux
    port map (
            O => \N__14275\,
            I => \N__14272\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__14272\,
            I => \Lab_UT.scctrl.g0_i_a7_2_0\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__14269\,
            I => \N__14266\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14263\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14260\
        );

    \I__2798\ : Span4Mux_v
    port map (
            O => \N__14260\,
            I => \N__14257\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__14257\,
            I => \Lab_UT.scctrl.next_state_1_i_a5_4_0_0\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14251\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__14251\,
            I => \Lab_UT.scctrl.N_8_0\
        );

    \I__2794\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14245\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__14245\,
            I => \Lab_UT.scctrl.g0_i_a9_1\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__14242\,
            I => \Lab_UT.scctrl.N_12_cascade_\
        );

    \I__2791\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14236\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__14236\,
            I => \Lab_UT.scctrl.g0_i_2\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__14233\,
            I => \N__14230\
        );

    \I__2788\ : InMux
    port map (
            O => \N__14230\,
            I => \N__14227\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__14227\,
            I => \N__14224\
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__14224\,
            I => \Lab_UT.scctrl.G_23_0_a9_0_0\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__14221\,
            I => \Lab_UT.scctrl.g0_i_a10_2_1_cascade_\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14215\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__14215\,
            I => \Lab_UT.scctrl.G_23_0_2\
        );

    \I__2782\ : InMux
    port map (
            O => \N__14212\,
            I => \N__14209\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__14209\,
            I => \Lab_UT.scctrl.N_2ctr\
        );

    \I__2780\ : InMux
    port map (
            O => \N__14206\,
            I => \N__14203\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__14203\,
            I => \Lab_UT.scctrl.g0_i_0\
        );

    \I__2778\ : InMux
    port map (
            O => \N__14200\,
            I => \N__14195\
        );

    \I__2777\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14189\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14198\,
            I => \N__14189\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__14195\,
            I => \N__14186\
        );

    \I__2774\ : InMux
    port map (
            O => \N__14194\,
            I => \N__14183\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__14189\,
            I => \Lab_UT.state_ret_13_RNIHUNI41_0\
        );

    \I__2772\ : Odrv4
    port map (
            O => \N__14186\,
            I => \Lab_UT.state_ret_13_RNIHUNI41_0\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__14183\,
            I => \Lab_UT.state_ret_13_RNIHUNI41_0\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__14176\,
            I => \Lab_UT.state_ret_13_RNIHUNI41_0_cascade_\
        );

    \I__2769\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14170\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__14170\,
            I => \N__14166\
        );

    \I__2767\ : InMux
    port map (
            O => \N__14169\,
            I => \N__14163\
        );

    \I__2766\ : Span4Mux_h
    port map (
            O => \N__14166\,
            I => \N__14160\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__14163\,
            I => \Lab_UT.scdp.key1_2\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__14160\,
            I => \Lab_UT.scdp.key1_2\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__14155\,
            I => \N__14150\
        );

    \I__2762\ : InMux
    port map (
            O => \N__14154\,
            I => \N__14147\
        );

    \I__2761\ : InMux
    port map (
            O => \N__14153\,
            I => \N__14141\
        );

    \I__2760\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14141\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__14147\,
            I => \N__14138\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14146\,
            I => \N__14135\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__14141\,
            I => \N__14132\
        );

    \I__2756\ : Span12Mux_s5_v
    port map (
            O => \N__14138\,
            I => \N__14129\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__14135\,
            I => \N__14124\
        );

    \I__2754\ : Span12Mux_s10_v
    port map (
            O => \N__14132\,
            I => \N__14124\
        );

    \I__2753\ : Odrv12
    port map (
            O => \N__14129\,
            I => \Lab_UT.sccDecrypt_0\
        );

    \I__2752\ : Odrv12
    port map (
            O => \N__14124\,
            I => \Lab_UT.sccDecrypt_0\
        );

    \I__2751\ : InMux
    port map (
            O => \N__14119\,
            I => \N__14114\
        );

    \I__2750\ : InMux
    port map (
            O => \N__14118\,
            I => \N__14109\
        );

    \I__2749\ : InMux
    port map (
            O => \N__14117\,
            I => \N__14109\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__14114\,
            I => \Lab_UT.state_ret_12_RNIMJCP8_0\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__14109\,
            I => \Lab_UT.state_ret_12_RNIMJCP8_0\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__14104\,
            I => \Lab_UT.sccDnibble2En_cascade_\
        );

    \I__2745\ : InMux
    port map (
            O => \N__14101\,
            I => \N__14098\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__14098\,
            I => \N__14095\
        );

    \I__2743\ : Span4Mux_h
    port map (
            O => \N__14095\,
            I => \N__14091\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14094\,
            I => \N__14088\
        );

    \I__2741\ : Span4Mux_v
    port map (
            O => \N__14091\,
            I => \N__14083\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__14088\,
            I => \N__14080\
        );

    \I__2739\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14077\
        );

    \I__2738\ : IoInMux
    port map (
            O => \N__14086\,
            I => \N__14074\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__14083\,
            I => \N__14069\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__14080\,
            I => \N__14069\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__14077\,
            I => \N__14066\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__14074\,
            I => \N__14063\
        );

    \I__2733\ : Span4Mux_h
    port map (
            O => \N__14069\,
            I => \N__14060\
        );

    \I__2732\ : Span4Mux_h
    port map (
            O => \N__14066\,
            I => \N__14057\
        );

    \I__2731\ : Span4Mux_s1_h
    port map (
            O => \N__14063\,
            I => \N__14054\
        );

    \I__2730\ : Odrv4
    port map (
            O => \N__14060\,
            I => \resetGen_rst_0_iso\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__14057\,
            I => \resetGen_rst_0_iso\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__14054\,
            I => \resetGen_rst_0_iso\
        );

    \I__2727\ : CEMux
    port map (
            O => \N__14047\,
            I => \N__14044\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__14044\,
            I => \Lab_UT.scdp.u1.sccDnibble2En_0\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14041\,
            I => \N__14037\
        );

    \I__2724\ : InMux
    port map (
            O => \N__14040\,
            I => \N__14034\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14037\,
            I => \N__14031\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__14034\,
            I => \N__14028\
        );

    \I__2721\ : Span4Mux_s2_v
    port map (
            O => \N__14031\,
            I => \N__14023\
        );

    \I__2720\ : Span4Mux_h
    port map (
            O => \N__14028\,
            I => \N__14023\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__14023\,
            I => \Lab_UT.scdp.N_37\
        );

    \I__2718\ : InMux
    port map (
            O => \N__14020\,
            I => \N__14014\
        );

    \I__2717\ : InMux
    port map (
            O => \N__14019\,
            I => \N__14014\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__14014\,
            I => \N__14010\
        );

    \I__2715\ : InMux
    port map (
            O => \N__14013\,
            I => \N__14007\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__14010\,
            I => \Lab_UT.sccDnibble2En\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__14007\,
            I => \Lab_UT.sccDnibble2En\
        );

    \I__2712\ : InMux
    port map (
            O => \N__14002\,
            I => \N__13998\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__14001\,
            I => \N__13995\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__13998\,
            I => \N__13992\
        );

    \I__2709\ : InMux
    port map (
            O => \N__13995\,
            I => \N__13989\
        );

    \I__2708\ : Span4Mux_h
    port map (
            O => \N__13992\,
            I => \N__13985\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__13989\,
            I => \N__13982\
        );

    \I__2706\ : InMux
    port map (
            O => \N__13988\,
            I => \N__13979\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__13985\,
            I => \N__13976\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__13982\,
            I => \N__13973\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__13979\,
            I => \Lab_UT.scdp.byteToDecrypt_1\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__13976\,
            I => \Lab_UT.scdp.byteToDecrypt_1\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__13973\,
            I => \Lab_UT.scdp.byteToDecrypt_1\
        );

    \I__2700\ : IoInMux
    port map (
            O => \N__13966\,
            I => \N__13960\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__13965\,
            I => \N__13957\
        );

    \I__2698\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13954\
        );

    \I__2697\ : InMux
    port map (
            O => \N__13963\,
            I => \N__13951\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__13960\,
            I => \N__13948\
        );

    \I__2695\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13945\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__13954\,
            I => \N__13942\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__13951\,
            I => \N__13939\
        );

    \I__2692\ : IoSpan4Mux
    port map (
            O => \N__13948\,
            I => \N__13936\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__13945\,
            I => \N__13933\
        );

    \I__2690\ : Span4Mux_v
    port map (
            O => \N__13942\,
            I => \N__13930\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__13939\,
            I => \N__13923\
        );

    \I__2688\ : Span4Mux_s1_v
    port map (
            O => \N__13936\,
            I => \N__13923\
        );

    \I__2687\ : Span4Mux_v
    port map (
            O => \N__13933\,
            I => \N__13923\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__13930\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__13923\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__13918\,
            I => \Lab_UT.scctrl.g0_i_a9_0_1_cascade_\
        );

    \I__2683\ : InMux
    port map (
            O => \N__13915\,
            I => \N__13912\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__13912\,
            I => \N__13908\
        );

    \I__2681\ : InMux
    port map (
            O => \N__13911\,
            I => \N__13905\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__13908\,
            I => \Lab_UT.scctrl.next_state77_2\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__13905\,
            I => \Lab_UT.scctrl.next_state77_2\
        );

    \I__2678\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13897\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__13897\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz_4\
        );

    \I__2676\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13891\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__13891\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__13888\,
            I => \N__13885\
        );

    \I__2673\ : InMux
    port map (
            O => \N__13885\,
            I => \N__13879\
        );

    \I__2672\ : InMux
    port map (
            O => \N__13884\,
            I => \N__13879\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__13879\,
            I => \N__13876\
        );

    \I__2670\ : Odrv12
    port map (
            O => \N__13876\,
            I => \Lab_UT.scctrl.next_state76\
        );

    \I__2669\ : InMux
    port map (
            O => \N__13873\,
            I => \N__13870\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__13870\,
            I => \N__13866\
        );

    \I__2667\ : InMux
    port map (
            O => \N__13869\,
            I => \N__13863\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__13866\,
            I => \N__13860\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__13863\,
            I => \Lab_UT.scdp.key2_3\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__13860\,
            I => \Lab_UT.scdp.key2_3\
        );

    \I__2663\ : InMux
    port map (
            O => \N__13855\,
            I => \N__13852\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__13852\,
            I => \N__13848\
        );

    \I__2661\ : InMux
    port map (
            O => \N__13851\,
            I => \N__13845\
        );

    \I__2660\ : Span4Mux_h
    port map (
            O => \N__13848\,
            I => \N__13842\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__13845\,
            I => \Lab_UT.scdp.key2_6\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__13842\,
            I => \Lab_UT.scdp.key2_6\
        );

    \I__2657\ : InMux
    port map (
            O => \N__13837\,
            I => \N__13831\
        );

    \I__2656\ : InMux
    port map (
            O => \N__13836\,
            I => \N__13828\
        );

    \I__2655\ : InMux
    port map (
            O => \N__13835\,
            I => \N__13823\
        );

    \I__2654\ : InMux
    port map (
            O => \N__13834\,
            I => \N__13823\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__13831\,
            I => \Lab_UT.state_ret_14_RNI416G41_0\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__13828\,
            I => \Lab_UT.state_ret_14_RNI416G41_0\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__13823\,
            I => \Lab_UT.state_ret_14_RNI416G41_0\
        );

    \I__2650\ : InMux
    port map (
            O => \N__13816\,
            I => \N__13812\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__13815\,
            I => \N__13809\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__13812\,
            I => \N__13806\
        );

    \I__2647\ : InMux
    port map (
            O => \N__13809\,
            I => \N__13803\
        );

    \I__2646\ : Span4Mux_h
    port map (
            O => \N__13806\,
            I => \N__13800\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__13803\,
            I => \Lab_UT.scdp.key3_6\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__13800\,
            I => \Lab_UT.scdp.key3_6\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__13795\,
            I => \N__13792\
        );

    \I__2642\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13788\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__13791\,
            I => \N__13785\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__13788\,
            I => \N__13782\
        );

    \I__2639\ : InMux
    port map (
            O => \N__13785\,
            I => \N__13779\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__13782\,
            I => \N__13776\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__13779\,
            I => \Lab_UT.scdp.key3_2\
        );

    \I__2636\ : Odrv4
    port map (
            O => \N__13776\,
            I => \Lab_UT.scdp.key3_2\
        );

    \I__2635\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13764\
        );

    \I__2634\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13759\
        );

    \I__2633\ : InMux
    port map (
            O => \N__13769\,
            I => \N__13759\
        );

    \I__2632\ : InMux
    port map (
            O => \N__13768\,
            I => \N__13754\
        );

    \I__2631\ : InMux
    port map (
            O => \N__13767\,
            I => \N__13754\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__13764\,
            I => \Lab_UT.state_2_RNI44QH41_0_2\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__13759\,
            I => \Lab_UT.state_2_RNI44QH41_0_2\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__13754\,
            I => \Lab_UT.state_2_RNI44QH41_0_2\
        );

    \I__2627\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13744\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__13744\,
            I => \N__13741\
        );

    \I__2625\ : Span4Mux_v
    port map (
            O => \N__13741\,
            I => \N__13737\
        );

    \I__2624\ : InMux
    port map (
            O => \N__13740\,
            I => \N__13734\
        );

    \I__2623\ : Span4Mux_s2_v
    port map (
            O => \N__13737\,
            I => \N__13731\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__13734\,
            I => \Lab_UT.scdp.key2_7\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__13731\,
            I => \Lab_UT.scdp.key2_7\
        );

    \I__2620\ : InMux
    port map (
            O => \N__13726\,
            I => \N__13719\
        );

    \I__2619\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13714\
        );

    \I__2618\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13714\
        );

    \I__2617\ : InMux
    port map (
            O => \N__13723\,
            I => \N__13711\
        );

    \I__2616\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13708\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__13719\,
            I => \Lab_UT.state_2_RNIF0RJ41_0_2\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__13714\,
            I => \Lab_UT.state_2_RNIF0RJ41_0_2\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__13711\,
            I => \Lab_UT.state_2_RNIF0RJ41_0_2\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__13708\,
            I => \Lab_UT.state_2_RNIF0RJ41_0_2\
        );

    \I__2611\ : InMux
    port map (
            O => \N__13699\,
            I => \N__13696\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__13696\,
            I => \N__13692\
        );

    \I__2609\ : InMux
    port map (
            O => \N__13695\,
            I => \N__13689\
        );

    \I__2608\ : Span4Mux_h
    port map (
            O => \N__13692\,
            I => \N__13686\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__13689\,
            I => \Lab_UT.scdp.key3_3\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__13686\,
            I => \Lab_UT.scdp.key3_3\
        );

    \I__2605\ : InMux
    port map (
            O => \N__13681\,
            I => \N__13677\
        );

    \I__2604\ : InMux
    port map (
            O => \N__13680\,
            I => \N__13674\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__13677\,
            I => \Lab_UT.scdp.key0_0\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__13674\,
            I => \Lab_UT.scdp.key0_0\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__13669\,
            I => \N__13666\
        );

    \I__2600\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13662\
        );

    \I__2599\ : InMux
    port map (
            O => \N__13665\,
            I => \N__13659\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__13662\,
            I => \Lab_UT.scdp.key0_2\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__13659\,
            I => \Lab_UT.scdp.key0_2\
        );

    \I__2596\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13650\
        );

    \I__2595\ : InMux
    port map (
            O => \N__13653\,
            I => \N__13647\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__13650\,
            I => \N__13644\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__13647\,
            I => \Lab_UT.scdp.key1_4\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__13644\,
            I => \Lab_UT.scdp.key1_4\
        );

    \I__2591\ : InMux
    port map (
            O => \N__13639\,
            I => \N__13632\
        );

    \I__2590\ : InMux
    port map (
            O => \N__13638\,
            I => \N__13629\
        );

    \I__2589\ : InMux
    port map (
            O => \N__13637\,
            I => \N__13626\
        );

    \I__2588\ : InMux
    port map (
            O => \N__13636\,
            I => \N__13621\
        );

    \I__2587\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13621\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__13632\,
            I => \N__13618\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__13629\,
            I => \Lab_UT.state_ret_13_RNIQ72741_0\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__13626\,
            I => \Lab_UT.state_ret_13_RNIQ72741_0\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__13621\,
            I => \Lab_UT.state_ret_13_RNIQ72741_0\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__13618\,
            I => \Lab_UT.state_ret_13_RNIQ72741_0\
        );

    \I__2581\ : InMux
    port map (
            O => \N__13609\,
            I => \N__13606\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__13606\,
            I => \N__13603\
        );

    \I__2579\ : Span4Mux_h
    port map (
            O => \N__13603\,
            I => \N__13599\
        );

    \I__2578\ : InMux
    port map (
            O => \N__13602\,
            I => \N__13596\
        );

    \I__2577\ : Span4Mux_h
    port map (
            O => \N__13599\,
            I => \N__13593\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__13596\,
            I => \Lab_UT.scdp.key1_6\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__13593\,
            I => \Lab_UT.scdp.key1_6\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__13588\,
            I => \Lab_UT.scctrl.next_state77_cascade_\
        );

    \I__2573\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13580\
        );

    \I__2572\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13575\
        );

    \I__2571\ : InMux
    port map (
            O => \N__13583\,
            I => \N__13575\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__13580\,
            I => \N__13572\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__13575\,
            I => \Lab_UT.scctrl.next_state_3_sqmuxa\
        );

    \I__2568\ : Odrv4
    port map (
            O => \N__13572\,
            I => \Lab_UT.scctrl.next_state_3_sqmuxa\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__13567\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_0_cascade_\
        );

    \I__2566\ : InMux
    port map (
            O => \N__13564\,
            I => \N__13561\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__13561\,
            I => \Lab_UT.scctrl.next_state77\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__13558\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_cascade_\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__13555\,
            I => \Lab_UT.scctrl.g0_i_a9_3_4_cascade_\
        );

    \I__2562\ : InMux
    port map (
            O => \N__13552\,
            I => \N__13549\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__13549\,
            I => \N__13546\
        );

    \I__2560\ : Span4Mux_s3_v
    port map (
            O => \N__13546\,
            I => \N__13543\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__13543\,
            I => \N__13540\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__13540\,
            I => \Lab_UT.scctrl.g0_i_a9_3_5\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__13537\,
            I => \Lab_UT.scctrl.next_state_1_0_a5_2_out_cascade_\
        );

    \I__2556\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13531\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__13531\,
            I => \Lab_UT.scctrl.N_222_1\
        );

    \I__2554\ : InMux
    port map (
            O => \N__13528\,
            I => \N__13525\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__13525\,
            I => \N__13522\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__13522\,
            I => \Lab_UT.scctrl.next_state_3_sqmuxa_0\
        );

    \I__2551\ : InMux
    port map (
            O => \N__13519\,
            I => \N__13516\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__13516\,
            I => \N__13513\
        );

    \I__2549\ : Odrv12
    port map (
            O => \N__13513\,
            I => \Lab_UT.scdp.a2b.g1_1_a3_0Z0Z_0\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__13510\,
            I => \N__13506\
        );

    \I__2547\ : InMux
    port map (
            O => \N__13509\,
            I => \N__13503\
        );

    \I__2546\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13500\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__13503\,
            I => \buart__rx_shifter_ret_1_fast\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__13500\,
            I => \buart__rx_shifter_ret_1_fast\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__13495\,
            I => \N__13492\
        );

    \I__2542\ : InMux
    port map (
            O => \N__13492\,
            I => \N__13489\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__13489\,
            I => \N__13486\
        );

    \I__2540\ : Odrv12
    port map (
            O => \N__13486\,
            I => \Lab_UT.scctrl.g0_i_o9_0Z0Z_2\
        );

    \I__2539\ : InMux
    port map (
            O => \N__13483\,
            I => \N__13477\
        );

    \I__2538\ : InMux
    port map (
            O => \N__13482\,
            I => \N__13477\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__13477\,
            I => \Lab_UT.dk.un4_de_hexZ0Z_1\
        );

    \I__2536\ : InMux
    port map (
            O => \N__13474\,
            I => \N__13470\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__13473\,
            I => \N__13465\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__13470\,
            I => \N__13461\
        );

    \I__2533\ : InMux
    port map (
            O => \N__13469\,
            I => \N__13456\
        );

    \I__2532\ : InMux
    port map (
            O => \N__13468\,
            I => \N__13456\
        );

    \I__2531\ : InMux
    port map (
            O => \N__13465\,
            I => \N__13453\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13450\
        );

    \I__2529\ : Span4Mux_h
    port map (
            O => \N__13461\,
            I => \N__13447\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__13456\,
            I => bu_rx_data_i_3_4
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__13453\,
            I => bu_rx_data_i_3_4
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13450\,
            I => bu_rx_data_i_3_4
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__13447\,
            I => bu_rx_data_i_3_4
        );

    \I__2524\ : InMux
    port map (
            O => \N__13438\,
            I => \N__13434\
        );

    \I__2523\ : InMux
    port map (
            O => \N__13437\,
            I => \N__13430\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__13434\,
            I => \N__13427\
        );

    \I__2521\ : InMux
    port map (
            O => \N__13433\,
            I => \N__13424\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__13430\,
            I => \N__13421\
        );

    \I__2519\ : Span4Mux_s3_h
    port map (
            O => \N__13427\,
            I => \N__13418\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__13424\,
            I => \N__13413\
        );

    \I__2517\ : Span4Mux_s3_h
    port map (
            O => \N__13421\,
            I => \N__13413\
        );

    \I__2516\ : Span4Mux_h
    port map (
            O => \N__13418\,
            I => \N__13401\
        );

    \I__2515\ : Span4Mux_h
    port map (
            O => \N__13413\,
            I => \N__13401\
        );

    \I__2514\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13396\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13411\,
            I => \N__13396\
        );

    \I__2512\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13385\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13409\,
            I => \N__13385\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13408\,
            I => \N__13385\
        );

    \I__2509\ : InMux
    port map (
            O => \N__13407\,
            I => \N__13385\
        );

    \I__2508\ : InMux
    port map (
            O => \N__13406\,
            I => \N__13385\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__13401\,
            I => bu_rx_data_5
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__13396\,
            I => bu_rx_data_5
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13385\,
            I => bu_rx_data_5
        );

    \I__2504\ : InMux
    port map (
            O => \N__13378\,
            I => \N__13370\
        );

    \I__2503\ : InMux
    port map (
            O => \N__13377\,
            I => \N__13365\
        );

    \I__2502\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13365\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13375\,
            I => \N__13358\
        );

    \I__2500\ : InMux
    port map (
            O => \N__13374\,
            I => \N__13358\
        );

    \I__2499\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13358\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__13370\,
            I => \N__13354\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__13365\,
            I => \N__13351\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__13358\,
            I => \N__13346\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13357\,
            I => \N__13343\
        );

    \I__2494\ : Span12Mux_s6_v
    port map (
            O => \N__13354\,
            I => \N__13338\
        );

    \I__2493\ : Span12Mux_s9_v
    port map (
            O => \N__13351\,
            I => \N__13338\
        );

    \I__2492\ : InMux
    port map (
            O => \N__13350\,
            I => \N__13333\
        );

    \I__2491\ : InMux
    port map (
            O => \N__13349\,
            I => \N__13333\
        );

    \I__2490\ : Odrv4
    port map (
            O => \N__13346\,
            I => bu_rx_data_4
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__13343\,
            I => bu_rx_data_4
        );

    \I__2488\ : Odrv12
    port map (
            O => \N__13338\,
            I => bu_rx_data_4
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__13333\,
            I => bu_rx_data_4
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__13324\,
            I => \N__13319\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__13323\,
            I => \N__13315\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__13322\,
            I => \N__13312\
        );

    \I__2483\ : InMux
    port map (
            O => \N__13319\,
            I => \N__13309\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13318\,
            I => \N__13306\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13315\,
            I => \N__13300\
        );

    \I__2480\ : InMux
    port map (
            O => \N__13312\,
            I => \N__13300\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__13309\,
            I => \N__13297\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__13306\,
            I => \N__13294\
        );

    \I__2477\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13291\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__13300\,
            I => \N__13288\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__13297\,
            I => bu_rx_data_i_2_6
        );

    \I__2474\ : Odrv12
    port map (
            O => \N__13294\,
            I => bu_rx_data_i_2_6
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__13291\,
            I => bu_rx_data_i_2_6
        );

    \I__2472\ : Odrv4
    port map (
            O => \N__13288\,
            I => bu_rx_data_i_2_6
        );

    \I__2471\ : InMux
    port map (
            O => \N__13279\,
            I => \N__13275\
        );

    \I__2470\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13272\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__13275\,
            I => \Lab_UT.un1_de_hex_2\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13272\,
            I => \Lab_UT.un1_de_hex_2\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__13267\,
            I => \Lab_UT.un1_de_hex_2_cascade_\
        );

    \I__2466\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13261\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__13261\,
            I => \Lab_UT.scctrl.N_9_0\
        );

    \I__2464\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13255\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__13255\,
            I => bu_rx_data_fast_0
        );

    \I__2462\ : InMux
    port map (
            O => \N__13252\,
            I => \N__13247\
        );

    \I__2461\ : InMux
    port map (
            O => \N__13251\,
            I => \N__13244\
        );

    \I__2460\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13241\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__13247\,
            I => \N__13238\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__13244\,
            I => \buart__rx_shifter_0_fast_3\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__13241\,
            I => \buart__rx_shifter_0_fast_3\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__13238\,
            I => \buart__rx_shifter_0_fast_3\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__13231\,
            I => \Lab_UT.dk.un7_de_hex_xZ0Z0_cascade_\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__13228\,
            I => \Lab_UT.dk.un7_de_hex_0_cascade_\
        );

    \I__2453\ : InMux
    port map (
            O => \N__13225\,
            I => \N__13222\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__13222\,
            I => \Lab_UT.dk.un7_de_hex_0\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__13219\,
            I => \Lab_UT.un4_de_hex_cascade_\
        );

    \I__2450\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13213\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13213\,
            I => \buart__rx_shifter_0_fast_1\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__13210\,
            I => \Lab_UT.scctrl.EmsLoaded_cascade_\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__13207\,
            I => \Lab_UT.sccElsBitsLd_cascade_\
        );

    \I__2446\ : CEMux
    port map (
            O => \N__13204\,
            I => \N__13201\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__13201\,
            I => \N__13197\
        );

    \I__2444\ : CEMux
    port map (
            O => \N__13200\,
            I => \N__13194\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__13197\,
            I => \N__13189\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__13194\,
            I => \N__13189\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__13189\,
            I => \N__13186\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__13186\,
            I => \Lab_UT.scdp.sccElsBitsLd_0\
        );

    \I__2439\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13174\
        );

    \I__2438\ : InMux
    port map (
            O => \N__13182\,
            I => \N__13174\
        );

    \I__2437\ : InMux
    port map (
            O => \N__13181\,
            I => \N__13174\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__13174\,
            I => \N__13171\
        );

    \I__2435\ : Span4Mux_v
    port map (
            O => \N__13171\,
            I => \N__13167\
        );

    \I__2434\ : InMux
    port map (
            O => \N__13170\,
            I => \N__13164\
        );

    \I__2433\ : Span4Mux_v
    port map (
            O => \N__13167\,
            I => \N__13161\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__13164\,
            I => \Lab_UT.sccElsBitsLd\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__13161\,
            I => \Lab_UT.sccElsBitsLd\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__13156\,
            I => \N__13153\
        );

    \I__2429\ : InMux
    port map (
            O => \N__13153\,
            I => \N__13150\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__13150\,
            I => \N__13147\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__13147\,
            I => \N__13143\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13146\,
            I => \N__13140\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__13143\,
            I => \Lab_UT.scdp.lsBitsi.lsBitsD_5\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__13140\,
            I => \Lab_UT.scdp.lsBitsi.lsBitsD_5\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__13135\,
            I => \Lab_UT_dk_de_cr_12_1_cascade_\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__13132\,
            I => \L4_PrintBuf_cascade_\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__13129\,
            I => \Lab_UT.sccDnibble1En_cascade_\
        );

    \I__2420\ : CEMux
    port map (
            O => \N__13126\,
            I => \N__13123\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__13123\,
            I => \N__13120\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__13120\,
            I => \N__13117\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__13117\,
            I => \Lab_UT.scdp.u0.sccDnibble1En_0\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__13114\,
            I => \Lab_UT.scctrl.next_state_1_sqmuxa_3_0_cascade_\
        );

    \I__2415\ : InMux
    port map (
            O => \N__13111\,
            I => \N__13105\
        );

    \I__2414\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13105\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__13105\,
            I => \N__13102\
        );

    \I__2412\ : Odrv4
    port map (
            O => \N__13102\,
            I => \Lab_UT.scctrl.state_retZ0Z_10\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__13099\,
            I => \Lab_UT.scctrl.next_state_1_sqmuxa_3_cascade_\
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__13096\,
            I => \N__13092\
        );

    \I__2409\ : InMux
    port map (
            O => \N__13095\,
            I => \N__13089\
        );

    \I__2408\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13086\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__13089\,
            I => \Lab_UT.scctrl.nibbleInZ0Z1\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13086\,
            I => \Lab_UT.scctrl.nibbleInZ0Z1\
        );

    \I__2405\ : CEMux
    port map (
            O => \N__13081\,
            I => \N__13078\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__13078\,
            I => \N__13075\
        );

    \I__2403\ : Span4Mux_v
    port map (
            O => \N__13075\,
            I => \N__13072\
        );

    \I__2402\ : Span4Mux_s2_v
    port map (
            O => \N__13072\,
            I => \N__13069\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__13069\,
            I => \Lab_UT.scctrl.N_1_0_i\
        );

    \I__2400\ : SRMux
    port map (
            O => \N__13066\,
            I => \N__13063\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__13063\,
            I => \N__13060\
        );

    \I__2398\ : Sp12to4
    port map (
            O => \N__13060\,
            I => \N__13056\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13053\
        );

    \I__2396\ : Odrv12
    port map (
            O => \N__13056\,
            I => \Lab_UT.scctrl.next_state_1_sqmuxa_3\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__13053\,
            I => \Lab_UT.scctrl.next_state_1_sqmuxa_3\
        );

    \I__2394\ : InMux
    port map (
            O => \N__13048\,
            I => \N__13045\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__13045\,
            I => \N__13041\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13044\,
            I => \N__13038\
        );

    \I__2391\ : Span12Mux_s3_v
    port map (
            O => \N__13041\,
            I => \N__13035\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__13038\,
            I => \Lab_UT.scctrl.un6_sccDecrypt\
        );

    \I__2389\ : Odrv12
    port map (
            O => \N__13035\,
            I => \Lab_UT.scctrl.un6_sccDecrypt\
        );

    \I__2388\ : InMux
    port map (
            O => \N__13030\,
            I => \N__13027\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__13027\,
            I => \N__13024\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__13024\,
            I => \Lab_UT.de_bigE\
        );

    \I__2385\ : InMux
    port map (
            O => \N__13021\,
            I => \N__13018\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__13018\,
            I => \N__13013\
        );

    \I__2383\ : InMux
    port map (
            O => \N__13017\,
            I => \N__13010\
        );

    \I__2382\ : InMux
    port map (
            O => \N__13016\,
            I => \N__13007\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__13013\,
            I => \Lab_UT.scctrl.next_state_1_i_a5_1_0\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__13010\,
            I => \Lab_UT.scctrl.next_state_1_i_a5_1_0\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__13007\,
            I => \Lab_UT.scctrl.next_state_1_i_a5_1_0\
        );

    \I__2378\ : InMux
    port map (
            O => \N__13000\,
            I => \N__12997\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__12997\,
            I => \Lab_UT.scctrl.EmsLoaded\
        );

    \I__2376\ : InMux
    port map (
            O => \N__12994\,
            I => \N__12991\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__12991\,
            I => \N__12988\
        );

    \I__2374\ : Odrv12
    port map (
            O => \N__12988\,
            I => \Lab_UT.scctrl.g0_7_1_0\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__12985\,
            I => \Lab_UT.scctrl.g2_0_2_cascade_\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__12982\,
            I => \Lab_UT.scctrl.g0_2_cascade_\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__12979\,
            I => \Lab_UT.scctrl.g0_7_cascade_\
        );

    \I__2370\ : InMux
    port map (
            O => \N__12976\,
            I => \N__12973\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__12973\,
            I => \Lab_UT.scctrl.g1_0\
        );

    \I__2368\ : InMux
    port map (
            O => \N__12970\,
            I => \N__12967\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__12967\,
            I => \N__12964\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__12964\,
            I => \Lab_UT.scctrl.g2_2\
        );

    \I__2365\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12958\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__12958\,
            I => \N__12955\
        );

    \I__2363\ : Odrv4
    port map (
            O => \N__12955\,
            I => \Lab_UT.scctrl.g1\
        );

    \I__2362\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12946\
        );

    \I__2361\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12946\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__12946\,
            I => \N__12942\
        );

    \I__2359\ : InMux
    port map (
            O => \N__12945\,
            I => \N__12939\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__12942\,
            I => \N__12936\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__12939\,
            I => \N__12933\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__12936\,
            I => \N__12930\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__12933\,
            I => \N__12927\
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__12930\,
            I => \Lab_UT.sccDnibble1En\
        );

    \I__2353\ : Odrv4
    port map (
            O => \N__12927\,
            I => \Lab_UT.sccDnibble1En\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__12922\,
            I => \Lab_UT.scctrl.next_state_rst_1_0_cascade_\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__12919\,
            I => \Lab_UT.scctrl.un1_state_3_1_reti_cascade_\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__12916\,
            I => \N__12913\
        );

    \I__2349\ : InMux
    port map (
            O => \N__12913\,
            I => \N__12910\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__12910\,
            I => \Lab_UT.de_bigE_0\
        );

    \I__2347\ : InMux
    port map (
            O => \N__12907\,
            I => \N__12903\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__12906\,
            I => \N__12900\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__12903\,
            I => \N__12897\
        );

    \I__2344\ : InMux
    port map (
            O => \N__12900\,
            I => \N__12894\
        );

    \I__2343\ : Span4Mux_h
    port map (
            O => \N__12897\,
            I => \N__12891\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__12894\,
            I => \Lab_UT.scdp.key3_1\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__12891\,
            I => \Lab_UT.scdp.key3_1\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__12886\,
            I => \N__12882\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__12885\,
            I => \N__12879\
        );

    \I__2338\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12876\
        );

    \I__2337\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12873\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__12876\,
            I => \N__12870\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__12873\,
            I => \Lab_UT.scdp.key1_0\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__12870\,
            I => \Lab_UT.scdp.key1_0\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__12865\,
            I => \N__12861\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__12864\,
            I => \N__12858\
        );

    \I__2331\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12855\
        );

    \I__2330\ : InMux
    port map (
            O => \N__12858\,
            I => \N__12852\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__12855\,
            I => \N__12849\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__12852\,
            I => \N__12846\
        );

    \I__2327\ : Odrv4
    port map (
            O => \N__12849\,
            I => \Lab_UT.scdp.key2_4\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__12846\,
            I => \Lab_UT.scdp.key2_4\
        );

    \I__2325\ : InMux
    port map (
            O => \N__12841\,
            I => \N__12838\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__12838\,
            I => \N__12834\
        );

    \I__2323\ : InMux
    port map (
            O => \N__12837\,
            I => \N__12831\
        );

    \I__2322\ : Span4Mux_h
    port map (
            O => \N__12834\,
            I => \N__12828\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__12831\,
            I => \Lab_UT.scdp.key3_4\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__12828\,
            I => \Lab_UT.scdp.key3_4\
        );

    \I__2319\ : InMux
    port map (
            O => \N__12823\,
            I => \N__12820\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__12820\,
            I => \N__12816\
        );

    \I__2317\ : InMux
    port map (
            O => \N__12819\,
            I => \N__12813\
        );

    \I__2316\ : Span4Mux_h
    port map (
            O => \N__12816\,
            I => \N__12810\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__12813\,
            I => \N__12807\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__12810\,
            I => \Lab_UT.sccEldByte\
        );

    \I__2313\ : Odrv12
    port map (
            O => \N__12807\,
            I => \Lab_UT.sccEldByte\
        );

    \I__2312\ : InMux
    port map (
            O => \N__12802\,
            I => \N__12769\
        );

    \I__2311\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12769\
        );

    \I__2310\ : InMux
    port map (
            O => \N__12800\,
            I => \N__12769\
        );

    \I__2309\ : InMux
    port map (
            O => \N__12799\,
            I => \N__12769\
        );

    \I__2308\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12769\
        );

    \I__2307\ : InMux
    port map (
            O => \N__12797\,
            I => \N__12769\
        );

    \I__2306\ : InMux
    port map (
            O => \N__12796\,
            I => \N__12769\
        );

    \I__2305\ : InMux
    port map (
            O => \N__12795\,
            I => \N__12769\
        );

    \I__2304\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12752\
        );

    \I__2303\ : InMux
    port map (
            O => \N__12793\,
            I => \N__12752\
        );

    \I__2302\ : InMux
    port map (
            O => \N__12792\,
            I => \N__12752\
        );

    \I__2301\ : InMux
    port map (
            O => \N__12791\,
            I => \N__12752\
        );

    \I__2300\ : InMux
    port map (
            O => \N__12790\,
            I => \N__12752\
        );

    \I__2299\ : InMux
    port map (
            O => \N__12789\,
            I => \N__12752\
        );

    \I__2298\ : InMux
    port map (
            O => \N__12788\,
            I => \N__12752\
        );

    \I__2297\ : InMux
    port map (
            O => \N__12787\,
            I => \N__12752\
        );

    \I__2296\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12733\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__12769\,
            I => \N__12728\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__12752\,
            I => \N__12728\
        );

    \I__2293\ : InMux
    port map (
            O => \N__12751\,
            I => \N__12713\
        );

    \I__2292\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12713\
        );

    \I__2291\ : InMux
    port map (
            O => \N__12749\,
            I => \N__12713\
        );

    \I__2290\ : InMux
    port map (
            O => \N__12748\,
            I => \N__12713\
        );

    \I__2289\ : InMux
    port map (
            O => \N__12747\,
            I => \N__12713\
        );

    \I__2288\ : InMux
    port map (
            O => \N__12746\,
            I => \N__12713\
        );

    \I__2287\ : InMux
    port map (
            O => \N__12745\,
            I => \N__12713\
        );

    \I__2286\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12710\
        );

    \I__2285\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12693\
        );

    \I__2284\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12693\
        );

    \I__2283\ : InMux
    port map (
            O => \N__12741\,
            I => \N__12693\
        );

    \I__2282\ : InMux
    port map (
            O => \N__12740\,
            I => \N__12693\
        );

    \I__2281\ : InMux
    port map (
            O => \N__12739\,
            I => \N__12693\
        );

    \I__2280\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12693\
        );

    \I__2279\ : InMux
    port map (
            O => \N__12737\,
            I => \N__12693\
        );

    \I__2278\ : InMux
    port map (
            O => \N__12736\,
            I => \N__12693\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__12733\,
            I => \N__12688\
        );

    \I__2276\ : Span4Mux_v
    port map (
            O => \N__12728\,
            I => \N__12688\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__12713\,
            I => \N__12683\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__12710\,
            I => \N__12683\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__12693\,
            I => \Lab_UT.state_ret_6_RNIL97G01_0\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__12688\,
            I => \Lab_UT.state_ret_6_RNIL97G01_0\
        );

    \I__2271\ : Odrv12
    port map (
            O => \N__12683\,
            I => \Lab_UT.state_ret_6_RNIL97G01_0\
        );

    \I__2270\ : IoInMux
    port map (
            O => \N__12676\,
            I => \N__12673\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__12673\,
            I => \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_iZ0\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__12670\,
            I => \Lab_UT.scctrl.un1_state_inv_cascade_\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__12667\,
            I => \Lab_UT.scctrl.state_ret_12_RNIUQFKZ0_cascade_\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__12664\,
            I => \Lab_UT.state_ret_12_RNIMJCP8_0_cascade_\
        );

    \I__2265\ : InMux
    port map (
            O => \N__12661\,
            I => \N__12658\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__12658\,
            I => \Lab_UT.scctrl.delayload\
        );

    \I__2263\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12651\
        );

    \I__2262\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12648\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__12651\,
            I => \N__12645\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__12648\,
            I => \N__12640\
        );

    \I__2259\ : Span4Mux_h
    port map (
            O => \N__12645\,
            I => \N__12640\
        );

    \I__2258\ : Span4Mux_v
    port map (
            O => \N__12640\,
            I => \N__12637\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__12637\,
            I => \Lab_UT.scctrl.delay3\
        );

    \I__2256\ : InMux
    port map (
            O => \N__12634\,
            I => \N__12631\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__12631\,
            I => \N__12628\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__12628\,
            I => \Lab_UT.scctrl.r4.delay4\
        );

    \I__2253\ : InMux
    port map (
            O => \N__12625\,
            I => \N__12622\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__12622\,
            I => \N__12619\
        );

    \I__2251\ : Span4Mux_v
    port map (
            O => \N__12619\,
            I => \N__12616\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__12616\,
            I => \Lab_UT.scdp.u1.byteToDecrypt_2\
        );

    \I__2249\ : InMux
    port map (
            O => \N__12613\,
            I => \N__12609\
        );

    \I__2248\ : InMux
    port map (
            O => \N__12612\,
            I => \N__12606\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12609\,
            I => \N__12603\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__12606\,
            I => \Lab_UT.scdp.key1_5\
        );

    \I__2245\ : Odrv12
    port map (
            O => \N__12603\,
            I => \Lab_UT.scdp.key1_5\
        );

    \I__2244\ : InMux
    port map (
            O => \N__12598\,
            I => \N__12594\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__12597\,
            I => \N__12591\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__12594\,
            I => \N__12588\
        );

    \I__2241\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12585\
        );

    \I__2240\ : Span4Mux_h
    port map (
            O => \N__12588\,
            I => \N__12582\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__12585\,
            I => \Lab_UT.scdp.key1_1\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__12582\,
            I => \Lab_UT.scdp.key1_1\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12577\,
            I => \N__12574\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__12574\,
            I => \N__12570\
        );

    \I__2235\ : InMux
    port map (
            O => \N__12573\,
            I => \N__12567\
        );

    \I__2234\ : Span12Mux_s5_h
    port map (
            O => \N__12570\,
            I => \N__12564\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__12567\,
            I => \Lab_UT.scdp.key2_5\
        );

    \I__2232\ : Odrv12
    port map (
            O => \N__12564\,
            I => \Lab_UT.scdp.key2_5\
        );

    \I__2231\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12555\
        );

    \I__2230\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12552\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__12555\,
            I => \N__12549\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__12552\,
            I => \Lab_UT.scdp.key3_5\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__12549\,
            I => \Lab_UT.scdp.key3_5\
        );

    \I__2226\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12541\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__12541\,
            I => \N__12537\
        );

    \I__2224\ : InMux
    port map (
            O => \N__12540\,
            I => \N__12534\
        );

    \I__2223\ : Span4Mux_h
    port map (
            O => \N__12537\,
            I => \N__12531\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__12534\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__12531\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0\
        );

    \I__2220\ : InMux
    port map (
            O => \N__12526\,
            I => \N__12523\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__12523\,
            I => \N__12519\
        );

    \I__2218\ : InMux
    port map (
            O => \N__12522\,
            I => \N__12516\
        );

    \I__2217\ : Span4Mux_h
    port map (
            O => \N__12519\,
            I => \N__12513\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__12516\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__12513\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12508\,
            I => \N__12504\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__12507\,
            I => \N__12501\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__12504\,
            I => \N__12497\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12492\
        );

    \I__2210\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12492\
        );

    \I__2209\ : Span4Mux_h
    port map (
            O => \N__12497\,
            I => \N__12489\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__12492\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_12\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__12489\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_12\
        );

    \I__2206\ : InMux
    port map (
            O => \N__12484\,
            I => \N__12480\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12483\,
            I => \N__12477\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__12480\,
            I => \N__12474\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__12477\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__12474\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13\
        );

    \I__2201\ : CEMux
    port map (
            O => \N__12469\,
            I => \N__12457\
        );

    \I__2200\ : CEMux
    port map (
            O => \N__12468\,
            I => \N__12457\
        );

    \I__2199\ : CEMux
    port map (
            O => \N__12467\,
            I => \N__12457\
        );

    \I__2198\ : CEMux
    port map (
            O => \N__12466\,
            I => \N__12457\
        );

    \I__2197\ : GlobalMux
    port map (
            O => \N__12457\,
            I => \N__12454\
        );

    \I__2196\ : gio2CtrlBuf
    port map (
            O => \N__12454\,
            I => \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_g\
        );

    \I__2195\ : InMux
    port map (
            O => \N__12451\,
            I => \N__12447\
        );

    \I__2194\ : InMux
    port map (
            O => \N__12450\,
            I => \N__12444\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__12447\,
            I => \Lab_UT.scdp.key3_0\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__12444\,
            I => \Lab_UT.scdp.key3_0\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12436\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__12436\,
            I => \N__12431\
        );

    \I__2189\ : InMux
    port map (
            O => \N__12435\,
            I => \N__12427\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__12434\,
            I => \N__12420\
        );

    \I__2187\ : Span4Mux_v
    port map (
            O => \N__12431\,
            I => \N__12416\
        );

    \I__2186\ : InMux
    port map (
            O => \N__12430\,
            I => \N__12413\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__12427\,
            I => \N__12410\
        );

    \I__2184\ : InMux
    port map (
            O => \N__12426\,
            I => \N__12405\
        );

    \I__2183\ : InMux
    port map (
            O => \N__12425\,
            I => \N__12405\
        );

    \I__2182\ : InMux
    port map (
            O => \N__12424\,
            I => \N__12400\
        );

    \I__2181\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12400\
        );

    \I__2180\ : InMux
    port map (
            O => \N__12420\,
            I => \N__12397\
        );

    \I__2179\ : InMux
    port map (
            O => \N__12419\,
            I => \N__12394\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__12416\,
            I => \buart__rx_bitcount_2\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__12413\,
            I => \buart__rx_bitcount_2\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__12410\,
            I => \buart__rx_bitcount_2\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__12405\,
            I => \buart__rx_bitcount_2\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__12400\,
            I => \buart__rx_bitcount_2\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__12397\,
            I => \buart__rx_bitcount_2\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__12394\,
            I => \buart__rx_bitcount_2\
        );

    \I__2171\ : InMux
    port map (
            O => \N__12379\,
            I => \N__12376\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12376\,
            I => \N__12373\
        );

    \I__2169\ : Span4Mux_v
    port map (
            O => \N__12373\,
            I => \N__12369\
        );

    \I__2168\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12366\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__12369\,
            I => \buart.Z_rx.bitcount_es_RNIGTPI1Z0Z_3\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__12366\,
            I => \buart.Z_rx.bitcount_es_RNIGTPI1Z0Z_3\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12361\,
            I => \N__12358\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__12358\,
            I => \N__12353\
        );

    \I__2163\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12348\
        );

    \I__2162\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12348\
        );

    \I__2161\ : Span4Mux_h
    port map (
            O => \N__12353\,
            I => \N__12345\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__12348\,
            I => \N__12342\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__12345\,
            I => \Lab_UT.scdp.d2eData_0\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__12342\,
            I => \Lab_UT.scdp.d2eData_0\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12334\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__12334\,
            I => \N__12330\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__12333\,
            I => \N__12327\
        );

    \I__2154\ : Span4Mux_v
    port map (
            O => \N__12330\,
            I => \N__12324\
        );

    \I__2153\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12321\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__12324\,
            I => \N__12318\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__12321\,
            I => \Lab_UT.scdp.lsBitsD_0\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__12318\,
            I => \Lab_UT.scdp.lsBitsD_0\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12309\
        );

    \I__2148\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12306\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__12309\,
            I => \N__12299\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__12306\,
            I => \N__12299\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12305\,
            I => \N__12294\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12304\,
            I => \N__12294\
        );

    \I__2143\ : Span4Mux_h
    port map (
            O => \N__12299\,
            I => \N__12291\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__12294\,
            I => \Lab_UT.scdp.lsBits_6\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__12291\,
            I => \Lab_UT.scdp.lsBits_6\
        );

    \I__2140\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12282\
        );

    \I__2139\ : InMux
    port map (
            O => \N__12285\,
            I => \N__12279\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__12282\,
            I => \N__12276\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__12279\,
            I => \N__12271\
        );

    \I__2136\ : Span4Mux_s3_v
    port map (
            O => \N__12276\,
            I => \N__12271\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__12271\,
            I => \Lab_UT.scdp.lsBitsD_4\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12268\,
            I => \N__12264\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__12267\,
            I => \N__12260\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__12264\,
            I => \N__12255\
        );

    \I__2131\ : InMux
    port map (
            O => \N__12263\,
            I => \N__12248\
        );

    \I__2130\ : InMux
    port map (
            O => \N__12260\,
            I => \N__12248\
        );

    \I__2129\ : InMux
    port map (
            O => \N__12259\,
            I => \N__12248\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12258\,
            I => \N__12245\
        );

    \I__2127\ : Span4Mux_h
    port map (
            O => \N__12255\,
            I => \N__12242\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__12248\,
            I => \N__12237\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__12245\,
            I => \N__12237\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__12242\,
            I => \N__12232\
        );

    \I__2123\ : Span4Mux_v
    port map (
            O => \N__12237\,
            I => \N__12232\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__12232\,
            I => \Lab_UT.scdp.N_48_i\
        );

    \I__2121\ : InMux
    port map (
            O => \N__12229\,
            I => \N__12226\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__12226\,
            I => \N__12223\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__12223\,
            I => \N__12220\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__12220\,
            I => \N__12216\
        );

    \I__2117\ : InMux
    port map (
            O => \N__12219\,
            I => \N__12213\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__12216\,
            I => \Lab_UT.scdp.N_52\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__12213\,
            I => \Lab_UT.scdp.N_52\
        );

    \I__2114\ : InMux
    port map (
            O => \N__12208\,
            I => \N__12204\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__12207\,
            I => \N__12201\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__12204\,
            I => \N__12198\
        );

    \I__2111\ : InMux
    port map (
            O => \N__12201\,
            I => \N__12195\
        );

    \I__2110\ : Span4Mux_h
    port map (
            O => \N__12198\,
            I => \N__12192\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__12195\,
            I => \N__12187\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__12192\,
            I => \N__12187\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__12187\,
            I => \Lab_UT.scdp.msBitsD_3\
        );

    \I__2106\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12181\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__12181\,
            I => \N__12172\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12169\
        );

    \I__2103\ : InMux
    port map (
            O => \N__12179\,
            I => \N__12166\
        );

    \I__2102\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12159\
        );

    \I__2101\ : InMux
    port map (
            O => \N__12177\,
            I => \N__12159\
        );

    \I__2100\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12159\
        );

    \I__2099\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12155\
        );

    \I__2098\ : Span4Mux_h
    port map (
            O => \N__12172\,
            I => \N__12152\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__12169\,
            I => \N__12149\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__12166\,
            I => \N__12146\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__12159\,
            I => \N__12143\
        );

    \I__2094\ : InMux
    port map (
            O => \N__12158\,
            I => \N__12140\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__12155\,
            I => \N__12137\
        );

    \I__2092\ : Span4Mux_v
    port map (
            O => \N__12152\,
            I => \N__12132\
        );

    \I__2091\ : Span4Mux_h
    port map (
            O => \N__12149\,
            I => \N__12132\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__12146\,
            I => \N__12127\
        );

    \I__2089\ : Span4Mux_v
    port map (
            O => \N__12143\,
            I => \N__12127\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__12140\,
            I => \N__12124\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__12137\,
            I => \buart__tx_uart_busy_0_i\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__12132\,
            I => \buart__tx_uart_busy_0_i\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__12127\,
            I => \buart__tx_uart_busy_0_i\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__12124\,
            I => \buart__tx_uart_busy_0_i\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__12115\,
            I => \N__12112\
        );

    \I__2082\ : InMux
    port map (
            O => \N__12112\,
            I => \N__12109\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__12109\,
            I => \N__12106\
        );

    \I__2080\ : Span4Mux_v
    port map (
            O => \N__12106\,
            I => \N__12100\
        );

    \I__2079\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12097\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__12104\,
            I => \N__12090\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__12103\,
            I => \N__12087\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__12100\,
            I => \N__12081\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__12097\,
            I => \N__12081\
        );

    \I__2074\ : InMux
    port map (
            O => \N__12096\,
            I => \N__12078\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12071\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12094\,
            I => \N__12071\
        );

    \I__2071\ : InMux
    port map (
            O => \N__12093\,
            I => \N__12071\
        );

    \I__2070\ : InMux
    port map (
            O => \N__12090\,
            I => \N__12064\
        );

    \I__2069\ : InMux
    port map (
            O => \N__12087\,
            I => \N__12064\
        );

    \I__2068\ : InMux
    port map (
            O => \N__12086\,
            I => \N__12064\
        );

    \I__2067\ : Span4Mux_v
    port map (
            O => \N__12081\,
            I => \N__12059\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__12078\,
            I => \N__12059\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__12071\,
            I => \buart.Z_tx.N_255\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__12064\,
            I => \buart.Z_tx.N_255\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__12059\,
            I => \buart.Z_tx.N_255\
        );

    \I__2062\ : InMux
    port map (
            O => \N__12052\,
            I => \N__12044\
        );

    \I__2061\ : InMux
    port map (
            O => \N__12051\,
            I => \N__12030\
        );

    \I__2060\ : InMux
    port map (
            O => \N__12050\,
            I => \N__12030\
        );

    \I__2059\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12025\
        );

    \I__2058\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12025\
        );

    \I__2057\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12022\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__12044\,
            I => \N__12019\
        );

    \I__2055\ : InMux
    port map (
            O => \N__12043\,
            I => \N__12012\
        );

    \I__2054\ : InMux
    port map (
            O => \N__12042\,
            I => \N__12012\
        );

    \I__2053\ : InMux
    port map (
            O => \N__12041\,
            I => \N__12012\
        );

    \I__2052\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12009\
        );

    \I__2051\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12002\
        );

    \I__2050\ : InMux
    port map (
            O => \N__12038\,
            I => \N__12002\
        );

    \I__2049\ : InMux
    port map (
            O => \N__12037\,
            I => \N__12002\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12036\,
            I => \N__11997\
        );

    \I__2047\ : InMux
    port map (
            O => \N__12035\,
            I => \N__11997\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__12030\,
            I => \N__11994\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__12025\,
            I => \N__11989\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__12022\,
            I => \N__11989\
        );

    \I__2043\ : Span12Mux_s9_v
    port map (
            O => \N__12019\,
            I => \N__11986\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__12012\,
            I => \N__11981\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__12009\,
            I => \N__11981\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__12002\,
            I => ufifo_utb_txdata_rdy_0
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__11997\,
            I => ufifo_utb_txdata_rdy_0
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__11994\,
            I => ufifo_utb_txdata_rdy_0
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__11989\,
            I => ufifo_utb_txdata_rdy_0
        );

    \I__2036\ : Odrv12
    port map (
            O => \N__11986\,
            I => ufifo_utb_txdata_rdy_0
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__11981\,
            I => ufifo_utb_txdata_rdy_0
        );

    \I__2034\ : InMux
    port map (
            O => \N__11968\,
            I => \N__11965\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__11965\,
            I => \N__11961\
        );

    \I__2032\ : InMux
    port map (
            O => \N__11964\,
            I => \N__11957\
        );

    \I__2031\ : Span4Mux_h
    port map (
            O => \N__11961\,
            I => \N__11954\
        );

    \I__2030\ : InMux
    port map (
            O => \N__11960\,
            I => \N__11951\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__11957\,
            I => \N__11948\
        );

    \I__2028\ : Span4Mux_v
    port map (
            O => \N__11954\,
            I => \N__11945\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__11951\,
            I => \N__11940\
        );

    \I__2026\ : Span12Mux_v
    port map (
            O => \N__11948\,
            I => \N__11940\
        );

    \I__2025\ : Odrv4
    port map (
            O => \N__11945\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__2024\ : Odrv12
    port map (
            O => \N__11940\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__2023\ : CascadeMux
    port map (
            O => \N__11935\,
            I => \N__11929\
        );

    \I__2022\ : InMux
    port map (
            O => \N__11934\,
            I => \N__11926\
        );

    \I__2021\ : InMux
    port map (
            O => \N__11933\,
            I => \N__11914\
        );

    \I__2020\ : InMux
    port map (
            O => \N__11932\,
            I => \N__11914\
        );

    \I__2019\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11914\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__11926\,
            I => \N__11911\
        );

    \I__2017\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11904\
        );

    \I__2016\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11904\
        );

    \I__2015\ : InMux
    port map (
            O => \N__11923\,
            I => \N__11904\
        );

    \I__2014\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11899\
        );

    \I__2013\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11899\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__11914\,
            I => \N__11894\
        );

    \I__2011\ : Span4Mux_v
    port map (
            O => \N__11911\,
            I => \N__11887\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__11904\,
            I => \N__11887\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__11899\,
            I => \N__11887\
        );

    \I__2008\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11882\
        );

    \I__2007\ : InMux
    port map (
            O => \N__11897\,
            I => \N__11882\
        );

    \I__2006\ : Span4Mux_v
    port map (
            O => \N__11894\,
            I => \N__11877\
        );

    \I__2005\ : Span4Mux_h
    port map (
            O => \N__11887\,
            I => \N__11877\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__11882\,
            I => bu_rx_data_3
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__11877\,
            I => bu_rx_data_3
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__11872\,
            I => \Lab_UT.scdp.a2b.N_53_cascade_\
        );

    \I__2001\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11866\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__11866\,
            I => \N__11862\
        );

    \I__1999\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11859\
        );

    \I__1998\ : Span4Mux_h
    port map (
            O => \N__11862\,
            I => \N__11856\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__11859\,
            I => \N__11851\
        );

    \I__1996\ : Span4Mux_v
    port map (
            O => \N__11856\,
            I => \N__11851\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__11851\,
            I => \Lab_UT.scdp.N_39\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__11848\,
            I => \N__11844\
        );

    \I__1993\ : InMux
    port map (
            O => \N__11847\,
            I => \N__11839\
        );

    \I__1992\ : InMux
    port map (
            O => \N__11844\,
            I => \N__11839\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__11839\,
            I => \N__11835\
        );

    \I__1990\ : InMux
    port map (
            O => \N__11838\,
            I => \N__11832\
        );

    \I__1989\ : Span4Mux_h
    port map (
            O => \N__11835\,
            I => \N__11829\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__11832\,
            I => \Lab_UT.scdp.byteToDecrypt_4\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__11829\,
            I => \Lab_UT.scdp.byteToDecrypt_4\
        );

    \I__1986\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11820\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__11823\,
            I => \N__11816\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__11820\,
            I => \N__11813\
        );

    \I__1983\ : InMux
    port map (
            O => \N__11819\,
            I => \N__11810\
        );

    \I__1982\ : InMux
    port map (
            O => \N__11816\,
            I => \N__11807\
        );

    \I__1981\ : Span4Mux_h
    port map (
            O => \N__11813\,
            I => \N__11804\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__11810\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_6\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__11807\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_6\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__11804\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_6\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__11797\,
            I => \N__11793\
        );

    \I__1976\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11790\
        );

    \I__1975\ : InMux
    port map (
            O => \N__11793\,
            I => \N__11787\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__11790\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__11787\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__11782\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsr_next_1_0_cascade_\
        );

    \I__1971\ : InMux
    port map (
            O => \N__11779\,
            I => \N__11774\
        );

    \I__1970\ : InMux
    port map (
            O => \N__11778\,
            I => \N__11771\
        );

    \I__1969\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11768\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__11774\,
            I => \N__11765\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__11771\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__11768\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__11765\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2\
        );

    \I__1964\ : InMux
    port map (
            O => \N__11758\,
            I => \N__11754\
        );

    \I__1963\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11751\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__11754\,
            I => \N__11748\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__11751\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_4\
        );

    \I__1960\ : Odrv4
    port map (
            O => \N__11748\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_4\
        );

    \I__1959\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11738\
        );

    \I__1958\ : InMux
    port map (
            O => \N__11742\,
            I => \N__11733\
        );

    \I__1957\ : InMux
    port map (
            O => \N__11741\,
            I => \N__11733\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__11738\,
            I => \N__11730\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__11733\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__11730\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5\
        );

    \I__1953\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11721\
        );

    \I__1952\ : InMux
    port map (
            O => \N__11724\,
            I => \N__11718\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__11721\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_11\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__11718\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_11\
        );

    \I__1949\ : InMux
    port map (
            O => \N__11713\,
            I => \N__11710\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__11710\,
            I => \Lab_UT.scctrl.next_state_0_sqmuxa_4Z0Z_0\
        );

    \I__1947\ : InMux
    port map (
            O => \N__11707\,
            I => \N__11704\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__11704\,
            I => \Lab_UT.dk.de_bigEZ0Z_1\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__11701\,
            I => \Lab_UT_dk_de_bigD_6_cascade_\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__11698\,
            I => \Lab_UT.de_bigE_cascade_\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__11695\,
            I => \Lab_UT.scdp.N_39_cascade_\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__11692\,
            I => \Lab_UT.scdp.a2b.N_50_cascade_\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__11689\,
            I => \N__11686\
        );

    \I__1940\ : InMux
    port map (
            O => \N__11686\,
            I => \N__11683\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__11683\,
            I => \Lab_UT.scdp.a2b.N_51\
        );

    \I__1938\ : InMux
    port map (
            O => \N__11680\,
            I => \N__11675\
        );

    \I__1937\ : InMux
    port map (
            O => \N__11679\,
            I => \N__11669\
        );

    \I__1936\ : InMux
    port map (
            O => \N__11678\,
            I => \N__11669\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__11675\,
            I => \N__11666\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__11674\,
            I => \N__11662\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__11669\,
            I => \N__11659\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__11666\,
            I => \N__11656\
        );

    \I__1931\ : InMux
    port map (
            O => \N__11665\,
            I => \N__11653\
        );

    \I__1930\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11650\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__11659\,
            I => bu_rx_data_i_2_5
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__11656\,
            I => bu_rx_data_i_2_5
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__11653\,
            I => bu_rx_data_i_2_5
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__11650\,
            I => bu_rx_data_i_2_5
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__11641\,
            I => \N__11638\
        );

    \I__1924\ : InMux
    port map (
            O => \N__11638\,
            I => \N__11635\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__11635\,
            I => \N__11632\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__11632\,
            I => \N__11629\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__11629\,
            I => \Lab_UT.scctrl.m24_e_5\
        );

    \I__1920\ : InMux
    port map (
            O => \N__11626\,
            I => \N__11623\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__11623\,
            I => \N__11620\
        );

    \I__1918\ : Span4Mux_v
    port map (
            O => \N__11620\,
            I => \N__11616\
        );

    \I__1917\ : InMux
    port map (
            O => \N__11619\,
            I => \N__11613\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__11616\,
            I => \Lab_UT.scdp.a2b.N_50\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__11613\,
            I => \Lab_UT.scdp.a2b.N_50\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__11608\,
            I => \bu_rx_data_rdy_cascade_\
        );

    \I__1913\ : InMux
    port map (
            O => \N__11605\,
            I => \N__11602\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__11602\,
            I => \Lab_UT.scctrl.delay1\
        );

    \I__1911\ : InMux
    port map (
            O => \N__11599\,
            I => \N__11596\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__11596\,
            I => \Lab_UT.scctrl.delay2\
        );

    \I__1909\ : InMux
    port map (
            O => \N__11593\,
            I => \N__11587\
        );

    \I__1908\ : InMux
    port map (
            O => \N__11592\,
            I => \N__11587\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__11587\,
            I => \N__11583\
        );

    \I__1906\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11580\
        );

    \I__1905\ : Span4Mux_v
    port map (
            O => \N__11583\,
            I => \N__11575\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__11580\,
            I => \N__11575\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__11575\,
            I => \N_6\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__11572\,
            I => \Lab_UT.scdp.pinst1.un12_pValidZ0Z_1_cascade_\
        );

    \I__1901\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11566\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__11566\,
            I => \Lab_UT.un7_pValid\
        );

    \I__1899\ : InMux
    port map (
            O => \N__11563\,
            I => \N__11557\
        );

    \I__1898\ : InMux
    port map (
            O => \N__11562\,
            I => \N__11557\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__11557\,
            I => \Lab_UT.un1_pValid\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__11554\,
            I => \Lab_UT.un7_pValid_cascade_\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__11551\,
            I => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_1_0_i_cascade_\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__11548\,
            I => \Lab_UT.g0_i_a9_1_3_cascade_\
        );

    \I__1893\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11542\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__11542\,
            I => \Lab_UT.scctrl.m24_e_4\
        );

    \I__1891\ : CascadeMux
    port map (
            O => \N__11539\,
            I => \Lab_UT.dk.escKey_4_reti_cascade_\
        );

    \I__1890\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11533\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__11533\,
            I => \N__11530\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__11530\,
            I => \Lab_UT.scctrl.g0_i_a7_1\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__11527\,
            I => \Lab_UT.scctrl.g0_i_a3_2_cascade_\
        );

    \I__1886\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11520\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__11523\,
            I => \N__11514\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__11520\,
            I => \N__11510\
        );

    \I__1883\ : InMux
    port map (
            O => \N__11519\,
            I => \N__11507\
        );

    \I__1882\ : InMux
    port map (
            O => \N__11518\,
            I => \N__11504\
        );

    \I__1881\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11501\
        );

    \I__1880\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11496\
        );

    \I__1879\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11496\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__11510\,
            I => \ufifo.tx_fsm.cstateZ0Z_4\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__11507\,
            I => \ufifo.tx_fsm.cstateZ0Z_4\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__11504\,
            I => \ufifo.tx_fsm.cstateZ0Z_4\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__11501\,
            I => \ufifo.tx_fsm.cstateZ0Z_4\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__11496\,
            I => \ufifo.tx_fsm.cstateZ0Z_4\
        );

    \I__1873\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11481\
        );

    \I__1872\ : InMux
    port map (
            O => \N__11484\,
            I => \N__11478\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__11481\,
            I => \ufifo.tx_fsm.N_59_0\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__11478\,
            I => \ufifo.tx_fsm.N_59_0\
        );

    \I__1869\ : InMux
    port map (
            O => \N__11473\,
            I => \N__11470\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__11470\,
            I => \N__11464\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11459\
        );

    \I__1866\ : InMux
    port map (
            O => \N__11468\,
            I => \N__11456\
        );

    \I__1865\ : InMux
    port map (
            O => \N__11467\,
            I => \N__11453\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__11464\,
            I => \N__11449\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11463\,
            I => \N__11444\
        );

    \I__1862\ : InMux
    port map (
            O => \N__11462\,
            I => \N__11444\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__11459\,
            I => \N__11439\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__11456\,
            I => \N__11436\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__11453\,
            I => \N__11433\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11452\,
            I => \N__11429\
        );

    \I__1857\ : Sp12to4
    port map (
            O => \N__11449\,
            I => \N__11424\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__11444\,
            I => \N__11424\
        );

    \I__1855\ : InMux
    port map (
            O => \N__11443\,
            I => \N__11419\
        );

    \I__1854\ : InMux
    port map (
            O => \N__11442\,
            I => \N__11419\
        );

    \I__1853\ : Span4Mux_h
    port map (
            O => \N__11439\,
            I => \N__11416\
        );

    \I__1852\ : Span4Mux_v
    port map (
            O => \N__11436\,
            I => \N__11411\
        );

    \I__1851\ : Span4Mux_h
    port map (
            O => \N__11433\,
            I => \N__11411\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11432\,
            I => \N__11408\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__11429\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1848\ : Odrv12
    port map (
            O => \N__11424\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__11419\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__11416\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__11411\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__11408\,
            I => \buart__tx_uart_busy_0\
        );

    \I__1843\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11391\
        );

    \I__1842\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11388\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__11391\,
            I => \N__11382\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__11388\,
            I => \N__11379\
        );

    \I__1839\ : InMux
    port map (
            O => \N__11387\,
            I => \N__11376\
        );

    \I__1838\ : InMux
    port map (
            O => \N__11386\,
            I => \N__11371\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__11385\,
            I => \N__11367\
        );

    \I__1836\ : Span4Mux_h
    port map (
            O => \N__11382\,
            I => \N__11364\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__11379\,
            I => \N__11359\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__11376\,
            I => \N__11359\
        );

    \I__1833\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11354\
        );

    \I__1832\ : InMux
    port map (
            O => \N__11374\,
            I => \N__11354\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__11371\,
            I => \N__11351\
        );

    \I__1830\ : InMux
    port map (
            O => \N__11370\,
            I => \N__11348\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11367\,
            I => \N__11345\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__11364\,
            I => \N__11340\
        );

    \I__1827\ : Span4Mux_h
    port map (
            O => \N__11359\,
            I => \N__11340\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__11354\,
            I => \N__11335\
        );

    \I__1825\ : Span12Mux_s11_v
    port map (
            O => \N__11351\,
            I => \N__11335\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__11348\,
            I => \ufifo.emitcrlf_fsm.cstateZ0Z_1\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__11345\,
            I => \ufifo.emitcrlf_fsm.cstateZ0Z_1\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__11340\,
            I => \ufifo.emitcrlf_fsm.cstateZ0Z_1\
        );

    \I__1821\ : Odrv12
    port map (
            O => \N__11335\,
            I => \ufifo.emitcrlf_fsm.cstateZ0Z_1\
        );

    \I__1820\ : InMux
    port map (
            O => \N__11326\,
            I => \N__11323\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__11323\,
            I => \ufifo.emitcrlf_fsm.cstate_srsts_rn_0_1\
        );

    \I__1818\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11316\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__11319\,
            I => \N__11313\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11316\,
            I => \N__11310\
        );

    \I__1815\ : InMux
    port map (
            O => \N__11313\,
            I => \N__11307\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__11310\,
            I => \ufifo.tx_fsm.cstateZ0Z_5\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__11307\,
            I => \ufifo.tx_fsm.cstateZ0Z_5\
        );

    \I__1812\ : InMux
    port map (
            O => \N__11302\,
            I => \N__11298\
        );

    \I__1811\ : InMux
    port map (
            O => \N__11301\,
            I => \N__11295\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__11298\,
            I => \N__11288\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__11295\,
            I => \N__11288\
        );

    \I__1808\ : InMux
    port map (
            O => \N__11294\,
            I => \N__11283\
        );

    \I__1807\ : InMux
    port map (
            O => \N__11293\,
            I => \N__11283\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__11288\,
            I => \N__11278\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__11283\,
            I => \N__11278\
        );

    \I__1804\ : Span4Mux_h
    port map (
            O => \N__11278\,
            I => \N__11275\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__11275\,
            I => \ufifo.crlfdone\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__11272\,
            I => \ufifo.tx_fsm.N_72_cascade_\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11257\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11268\,
            I => \N__11257\
        );

    \I__1799\ : InMux
    port map (
            O => \N__11267\,
            I => \N__11246\
        );

    \I__1798\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11246\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11246\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11246\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11263\,
            I => \N__11246\
        );

    \I__1794\ : InMux
    port map (
            O => \N__11262\,
            I => \N__11243\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__11257\,
            I => \N__11238\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__11246\,
            I => \N__11233\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__11243\,
            I => \N__11233\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11230\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11227\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__11238\,
            I => \N__11218\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__11233\,
            I => \N__11218\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__11230\,
            I => \N__11218\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__11227\,
            I => \N__11215\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11210\
        );

    \I__1783\ : InMux
    port map (
            O => \N__11225\,
            I => \N__11210\
        );

    \I__1782\ : Span4Mux_h
    port map (
            O => \N__11218\,
            I => \N__11207\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__11215\,
            I => \ufifo.cstate_0\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11210\,
            I => \ufifo.cstate_0\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__11207\,
            I => \ufifo.cstate_0\
        );

    \I__1778\ : InMux
    port map (
            O => \N__11200\,
            I => \N__11197\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__11197\,
            I => \Lab_UT.dk.de_bigEZ0Z_2\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__11194\,
            I => \Lab_UT.scdp.d2eData_3_5_cascade_\
        );

    \I__1775\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11188\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__11188\,
            I => \N__11185\
        );

    \I__1773\ : Span4Mux_h
    port map (
            O => \N__11185\,
            I => \N__11180\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11184\,
            I => \N__11175\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11175\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__11180\,
            I => \Lab_UT.scdp.e2dData_5\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__11175\,
            I => \Lab_UT.scdp.e2dData_5\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11164\
        );

    \I__1767\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11164\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__11164\,
            I => \Lab_UT.scdp.u0.byteToDecrypt_5\
        );

    \I__1765\ : InMux
    port map (
            O => \N__11161\,
            I => \N__11157\
        );

    \I__1764\ : InMux
    port map (
            O => \N__11160\,
            I => \N__11154\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__11157\,
            I => \Lab_UT.scdp.u0.byteToDecrypt_7\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__11154\,
            I => \Lab_UT.scdp.u0.byteToDecrypt_7\
        );

    \I__1761\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11144\
        );

    \I__1760\ : InMux
    port map (
            O => \N__11148\,
            I => \N__11141\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11138\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__11144\,
            I => \N__11131\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__11141\,
            I => \N__11131\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__11138\,
            I => \N__11131\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__11131\,
            I => \N__11128\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__11128\,
            I => \Lab_UT.scdp.val_0_3\
        );

    \I__1753\ : InMux
    port map (
            O => \N__11125\,
            I => \N__11122\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__11122\,
            I => \N__11118\
        );

    \I__1751\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11115\
        );

    \I__1750\ : Span4Mux_h
    port map (
            O => \N__11118\,
            I => \N__11112\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__11115\,
            I => \Lab_UT.scdp.key1_7\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__11112\,
            I => \Lab_UT.scdp.key1_7\
        );

    \I__1747\ : InMux
    port map (
            O => \N__11107\,
            I => \N__11103\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11106\,
            I => \N__11100\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__11103\,
            I => \N__11097\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__11100\,
            I => \Lab_UT.scdp.key1_3\
        );

    \I__1743\ : Odrv12
    port map (
            O => \N__11097\,
            I => \Lab_UT.scdp.key1_3\
        );

    \I__1742\ : SRMux
    port map (
            O => \N__11092\,
            I => \N__11087\
        );

    \I__1741\ : CEMux
    port map (
            O => \N__11091\,
            I => \N__11084\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__11090\,
            I => \N__11080\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__11087\,
            I => \N__11077\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__11084\,
            I => \N__11074\
        );

    \I__1737\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11071\
        );

    \I__1736\ : InMux
    port map (
            O => \N__11080\,
            I => \N__11068\
        );

    \I__1735\ : Span4Mux_h
    port map (
            O => \N__11077\,
            I => \N__11063\
        );

    \I__1734\ : Span4Mux_h
    port map (
            O => \N__11074\,
            I => \N__11063\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__11071\,
            I => \N__11058\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__11068\,
            I => \N__11058\
        );

    \I__1731\ : Sp12to4
    port map (
            O => \N__11063\,
            I => \N__11053\
        );

    \I__1730\ : Span12Mux_s4_h
    port map (
            O => \N__11058\,
            I => \N__11053\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__11053\,
            I => \ufifo.txDataValidDZ0\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11050\,
            I => \N__11047\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__11047\,
            I => \ufifo.emitcrlf_fsm.cstate_srsts_sn_1\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__11044\,
            I => \ufifo.N_57_0_1_cascade_\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11036\
        );

    \I__1724\ : InMux
    port map (
            O => \N__11040\,
            I => \N__11033\
        );

    \I__1723\ : InMux
    port map (
            O => \N__11039\,
            I => \N__11030\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__11036\,
            I => \N__11027\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__11033\,
            I => \N__11024\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__11030\,
            I => \N__11017\
        );

    \I__1719\ : Span4Mux_h
    port map (
            O => \N__11027\,
            I => \N__11017\
        );

    \I__1718\ : Span4Mux_h
    port map (
            O => \N__11024\,
            I => \N__11017\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__11017\,
            I => \Lab_UT.scdp.prng_lfsr_23\
        );

    \I__1716\ : InMux
    port map (
            O => \N__11014\,
            I => \N__11010\
        );

    \I__1715\ : CascadeMux
    port map (
            O => \N__11013\,
            I => \N__11007\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__11010\,
            I => \N__11004\
        );

    \I__1713\ : InMux
    port map (
            O => \N__11007\,
            I => \N__11001\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__11004\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__11001\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24\
        );

    \I__1710\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10992\
        );

    \I__1709\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10989\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__10992\,
            I => \N__10986\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__10989\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__10986\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19\
        );

    \I__1705\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10977\
        );

    \I__1704\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10974\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__10977\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__10974\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__10969\,
            I => \N__10965\
        );

    \I__1700\ : InMux
    port map (
            O => \N__10968\,
            I => \N__10962\
        );

    \I__1699\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10959\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__10962\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__10959\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28\
        );

    \I__1696\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10951\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__10951\,
            I => \N__10946\
        );

    \I__1694\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10943\
        );

    \I__1693\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10940\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__10946\,
            I => \N__10937\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__10943\,
            I => \N__10932\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__10940\,
            I => \N__10932\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__10937\,
            I => \Lab_UT.scdp.prng_lfsr_7\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__10932\,
            I => \Lab_UT.scdp.prng_lfsr_7\
        );

    \I__1687\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10923\
        );

    \I__1686\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10920\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__10923\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__10920\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__10915\,
            I => \N__10911\
        );

    \I__1682\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10908\
        );

    \I__1681\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10905\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__10908\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__10905\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__10900\,
            I => \N__10896\
        );

    \I__1677\ : InMux
    port map (
            O => \N__10899\,
            I => \N__10893\
        );

    \I__1676\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10890\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__10893\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__10890\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27\
        );

    \I__1673\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10881\
        );

    \I__1672\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10878\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__10881\,
            I => \N__10875\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__10878\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__10875\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21\
        );

    \I__1668\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10866\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__10869\,
            I => \N__10863\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__10866\,
            I => \N__10860\
        );

    \I__1665\ : InMux
    port map (
            O => \N__10863\,
            I => \N__10857\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__10860\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__10857\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29\
        );

    \I__1662\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10849\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__10849\,
            I => \N__10846\
        );

    \I__1660\ : Span4Mux_v
    port map (
            O => \N__10846\,
            I => \N__10843\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__10843\,
            I => \Lab_UT.scdp.d2eData_3_5\
        );

    \I__1658\ : InMux
    port map (
            O => \N__10840\,
            I => \N__10836\
        );

    \I__1657\ : InMux
    port map (
            O => \N__10839\,
            I => \N__10833\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__10836\,
            I => \N__10830\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__10833\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__10830\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22\
        );

    \I__1653\ : InMux
    port map (
            O => \N__10825\,
            I => \N__10821\
        );

    \I__1652\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10818\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__10821\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__10818\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__10813\,
            I => \N__10809\
        );

    \I__1648\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10806\
        );

    \I__1647\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10803\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__10806\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__10803\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25\
        );

    \I__1644\ : InMux
    port map (
            O => \N__10798\,
            I => \N__10794\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__10797\,
            I => \N__10791\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__10794\,
            I => \N__10787\
        );

    \I__1641\ : InMux
    port map (
            O => \N__10791\,
            I => \N__10784\
        );

    \I__1640\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10781\
        );

    \I__1639\ : Span4Mux_h
    port map (
            O => \N__10787\,
            I => \N__10778\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__10784\,
            I => \N__10775\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__10781\,
            I => \Lab_UT.scdp.prng_lfsr_15\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__10778\,
            I => \Lab_UT.scdp.prng_lfsr_15\
        );

    \I__1635\ : Odrv4
    port map (
            O => \N__10775\,
            I => \Lab_UT.scdp.prng_lfsr_15\
        );

    \I__1634\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10764\
        );

    \I__1633\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10761\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__10764\,
            I => \N__10758\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__10761\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__10758\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16\
        );

    \I__1629\ : InMux
    port map (
            O => \N__10753\,
            I => \N__10749\
        );

    \I__1628\ : InMux
    port map (
            O => \N__10752\,
            I => \N__10746\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__10749\,
            I => \N__10743\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__10746\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_3\
        );

    \I__1625\ : Odrv4
    port map (
            O => \N__10743\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_3\
        );

    \I__1624\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10734\
        );

    \I__1623\ : InMux
    port map (
            O => \N__10737\,
            I => \N__10731\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__10734\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__10731\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9\
        );

    \I__1620\ : InMux
    port map (
            O => \N__10726\,
            I => \N__10722\
        );

    \I__1619\ : InMux
    port map (
            O => \N__10725\,
            I => \N__10719\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__10722\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__10719\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10\
        );

    \I__1616\ : InMux
    port map (
            O => \N__10714\,
            I => \N__10711\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__10711\,
            I => \N__10707\
        );

    \I__1614\ : InMux
    port map (
            O => \N__10710\,
            I => \N__10704\
        );

    \I__1613\ : Span4Mux_h
    port map (
            O => \N__10707\,
            I => \N__10701\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__10704\,
            I => \N__10698\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__10701\,
            I => \N__10695\
        );

    \I__1610\ : Odrv12
    port map (
            O => \N__10698\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__10695\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__1608\ : InMux
    port map (
            O => \N__10690\,
            I => \N__10686\
        );

    \I__1607\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10683\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__10686\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__10683\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17\
        );

    \I__1604\ : InMux
    port map (
            O => \N__10678\,
            I => \N__10674\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10677\,
            I => \N__10671\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__10674\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_14\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__10671\,
            I => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_14\
        );

    \I__1600\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10660\
        );

    \I__1599\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10660\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__10660\,
            I => \Lab_UT.de_bigL_0\
        );

    \I__1597\ : InMux
    port map (
            O => \N__10657\,
            I => \N__10653\
        );

    \I__1596\ : InMux
    port map (
            O => \N__10656\,
            I => \N__10644\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__10653\,
            I => \N__10641\
        );

    \I__1594\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10636\
        );

    \I__1593\ : InMux
    port map (
            O => \N__10651\,
            I => \N__10636\
        );

    \I__1592\ : InMux
    port map (
            O => \N__10650\,
            I => \N__10633\
        );

    \I__1591\ : InMux
    port map (
            O => \N__10649\,
            I => \N__10630\
        );

    \I__1590\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10627\
        );

    \I__1589\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10624\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__10644\,
            I => \buart__rx_bitcount_3\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__10641\,
            I => \buart__rx_bitcount_3\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__10636\,
            I => \buart__rx_bitcount_3\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__10633\,
            I => \buart__rx_bitcount_3\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__10630\,
            I => \buart__rx_bitcount_3\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__10627\,
            I => \buart__rx_bitcount_3\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__10624\,
            I => \buart__rx_bitcount_3\
        );

    \I__1581\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10605\
        );

    \I__1580\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10600\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__10605\,
            I => \N__10595\
        );

    \I__1578\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10592\
        );

    \I__1577\ : InMux
    port map (
            O => \N__10603\,
            I => \N__10586\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__10600\,
            I => \N__10583\
        );

    \I__1575\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10578\
        );

    \I__1574\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10578\
        );

    \I__1573\ : Span4Mux_h
    port map (
            O => \N__10595\,
            I => \N__10573\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__10592\,
            I => \N__10573\
        );

    \I__1571\ : InMux
    port map (
            O => \N__10591\,
            I => \N__10570\
        );

    \I__1570\ : InMux
    port map (
            O => \N__10590\,
            I => \N__10565\
        );

    \I__1569\ : InMux
    port map (
            O => \N__10589\,
            I => \N__10565\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__10586\,
            I => \buart__rx_bitcount_0\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__10583\,
            I => \buart__rx_bitcount_0\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__10578\,
            I => \buart__rx_bitcount_0\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__10573\,
            I => \buart__rx_bitcount_0\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__10570\,
            I => \buart__rx_bitcount_0\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__10565\,
            I => \buart__rx_bitcount_0\
        );

    \I__1562\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10541\
        );

    \I__1561\ : InMux
    port map (
            O => \N__10551\,
            I => \N__10541\
        );

    \I__1560\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10536\
        );

    \I__1559\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10536\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__10548\,
            I => \N__10531\
        );

    \I__1557\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10528\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10525\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__10541\,
            I => \N__10522\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__10536\,
            I => \N__10519\
        );

    \I__1553\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10516\
        );

    \I__1552\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10511\
        );

    \I__1551\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10511\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__10528\,
            I => \buart__rx_bitcount_1\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__10525\,
            I => \buart__rx_bitcount_1\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__10522\,
            I => \buart__rx_bitcount_1\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__10519\,
            I => \buart__rx_bitcount_1\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__10516\,
            I => \buart__rx_bitcount_1\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__10511\,
            I => \buart__rx_bitcount_1\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__10498\,
            I => \N__10491\
        );

    \I__1543\ : InMux
    port map (
            O => \N__10497\,
            I => \N__10487\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10496\,
            I => \N__10481\
        );

    \I__1541\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10481\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10494\,
            I => \N__10478\
        );

    \I__1539\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10474\
        );

    \I__1538\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10471\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__10487\,
            I => \N__10468\
        );

    \I__1536\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10465\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__10481\,
            I => \N__10460\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__10478\,
            I => \N__10460\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10457\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__10474\,
            I => \buart__rx_bitcount_4\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__10471\,
            I => \buart__rx_bitcount_4\
        );

    \I__1530\ : Odrv12
    port map (
            O => \N__10468\,
            I => \buart__rx_bitcount_4\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__10465\,
            I => \buart__rx_bitcount_4\
        );

    \I__1528\ : Odrv4
    port map (
            O => \N__10460\,
            I => \buart__rx_bitcount_4\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__10457\,
            I => \buart__rx_bitcount_4\
        );

    \I__1526\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10441\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__10441\,
            I => \buart.Z_rx.shifter_0_fast_RNI1CIH1Z0Z_2\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__10438\,
            I => \buart.Z_rx.bitcount_es_RNIF6D61Z0Z_4_cascade_\
        );

    \I__1523\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10432\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__10432\,
            I => \Lab_UT_dk_de_bigD_0\
        );

    \I__1521\ : InMux
    port map (
            O => \N__10429\,
            I => \N__10426\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__10426\,
            I => \Lab_UT.dk.de_bigD_sxZ0\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__10423\,
            I => \Lab_UT_dk_de_bigD_0_cascade_\
        );

    \I__1518\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10416\
        );

    \I__1517\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10413\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__10416\,
            I => \Lab_UT.dk.de_bigD_1Z0Z_0\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__10413\,
            I => \Lab_UT.dk.de_bigD_1Z0Z_0\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__10408\,
            I => \N__10405\
        );

    \I__1513\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10402\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__10402\,
            I => \N__10399\
        );

    \I__1511\ : Span4Mux_h
    port map (
            O => \N__10399\,
            I => \N__10396\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__10396\,
            I => \buart.Z_rx.N_41_i_1\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__10393\,
            I => \N__10390\
        );

    \I__1508\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10387\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__10387\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10384\,
            I => \N__10381\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__10381\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__10378\,
            I => \N__10374\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10377\,
            I => \N__10368\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10374\,
            I => \N__10368\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__10373\,
            I => \N__10361\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__10368\,
            I => \N__10354\
        );

    \I__1499\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10351\
        );

    \I__1498\ : InMux
    port map (
            O => \N__10366\,
            I => \N__10346\
        );

    \I__1497\ : InMux
    port map (
            O => \N__10365\,
            I => \N__10346\
        );

    \I__1496\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10343\
        );

    \I__1495\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10334\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10360\,
            I => \N__10334\
        );

    \I__1493\ : InMux
    port map (
            O => \N__10359\,
            I => \N__10334\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10334\
        );

    \I__1491\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10331\
        );

    \I__1490\ : Span4Mux_v
    port map (
            O => \N__10354\,
            I => \N__10328\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__10351\,
            I => \N__10321\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__10346\,
            I => \N__10321\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__10343\,
            I => \N__10321\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__10334\,
            I => \N__10314\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__10331\,
            I => \N__10314\
        );

    \I__1484\ : Span4Mux_h
    port map (
            O => \N__10328\,
            I => \N__10314\
        );

    \I__1483\ : Odrv12
    port map (
            O => \N__10321\,
            I => \buart.Z_rx.startbit\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__10314\,
            I => \buart.Z_rx.startbit\
        );

    \I__1481\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10296\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10308\,
            I => \N__10296\
        );

    \I__1479\ : InMux
    port map (
            O => \N__10307\,
            I => \N__10296\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10296\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10293\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__10296\,
            I => \buart.Z_rx.N_45\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__10293\,
            I => \buart.Z_rx.N_45\
        );

    \I__1474\ : CascadeMux
    port map (
            O => \N__10288\,
            I => \N__10285\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10285\,
            I => \N__10282\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10282\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__1471\ : CEMux
    port map (
            O => \N__10279\,
            I => \N__10275\
        );

    \I__1470\ : CEMux
    port map (
            O => \N__10278\,
            I => \N__10272\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__10275\,
            I => \N__10269\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__10272\,
            I => \N__10266\
        );

    \I__1467\ : Span4Mux_v
    port map (
            O => \N__10269\,
            I => \N__10263\
        );

    \I__1466\ : Odrv4
    port map (
            O => \N__10266\,
            I => \buart.Z_rx.N_43\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__10263\,
            I => \buart.Z_rx.N_43\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__10258\,
            I => \N__10255\
        );

    \I__1463\ : InMux
    port map (
            O => \N__10255\,
            I => \N__10252\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__10252\,
            I => \Lab_UT.dk.de_bigL_sxZ0\
        );

    \I__1461\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10246\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__10246\,
            I => \Lab_UT.de_bigL_3\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10240\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__10240\,
            I => \N__10237\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__10237\,
            I => \Lab_UT.scctrl.g0_17_N_3LZ0Z3\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__10234\,
            I => \Lab_UT.de_bigL_3_cascade_\
        );

    \I__1455\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10228\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__10228\,
            I => \N__10225\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__10225\,
            I => \Lab_UT.scctrl.g0_17_N_2LZ0Z1\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__10222\,
            I => \buart.Z_rx.N_58_cascade_\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10219\,
            I => \N__10216\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__10216\,
            I => \N__10213\
        );

    \I__1449\ : Span4Mux_h
    port map (
            O => \N__10213\,
            I => \N__10209\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10212\,
            I => \N__10206\
        );

    \I__1447\ : Span4Mux_v
    port map (
            O => \N__10209\,
            I => \N__10203\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__10206\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__10203\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10194\
        );

    \I__1443\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10191\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__10194\,
            I => \buart.Z_rx.N_58\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__10191\,
            I => \buart.Z_rx.N_58\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__10186\,
            I => \buart.Z_rx.startbit_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10179\
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__10182\,
            I => \N__10175\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__10179\,
            I => \N__10172\
        );

    \I__1436\ : InMux
    port map (
            O => \N__10178\,
            I => \N__10167\
        );

    \I__1435\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10164\
        );

    \I__1434\ : Span4Mux_h
    port map (
            O => \N__10172\,
            I => \N__10161\
        );

    \I__1433\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10156\
        );

    \I__1432\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10156\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__10167\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__10164\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__10161\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__10156\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1427\ : InMux
    port map (
            O => \N__10147\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10144\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10141\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__1424\ : InMux
    port map (
            O => \N__10138\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__10135\,
            I => \N__10131\
        );

    \I__1422\ : InMux
    port map (
            O => \N__10134\,
            I => \N__10128\
        );

    \I__1421\ : InMux
    port map (
            O => \N__10131\,
            I => \N__10125\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10128\,
            I => \N__10122\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__10125\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__1418\ : Odrv4
    port map (
            O => \N__10122\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__10117\,
            I => \N__10113\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10116\,
            I => \N__10110\
        );

    \I__1415\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10107\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__10110\,
            I => \N__10104\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__10107\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__10104\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1411\ : CascadeMux
    port map (
            O => \N__10099\,
            I => \N__10096\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10096\,
            I => \N__10092\
        );

    \I__1409\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10089\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__10092\,
            I => \N__10086\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__10089\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1406\ : Odrv12
    port map (
            O => \N__10086\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1405\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10078\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__10078\,
            I => \ufifo.fifo.un1_emptyB_NE_2\
        );

    \I__1403\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10072\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__10072\,
            I => \N__10069\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__10069\,
            I => \ufifo.fifo.un1_emptyB_NE_1\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__10066\,
            I => \N__10063\
        );

    \I__1399\ : InMux
    port map (
            O => \N__10063\,
            I => \N__10060\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__10060\,
            I => \N__10057\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__10057\,
            I => \ufifo.fifo.un1_emptyB_NE_3\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10054\,
            I => \N__10051\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__10051\,
            I => \N__10048\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__10048\,
            I => \ufifo.fifo.un1_emptyB_NE_4\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__10045\,
            I => \ufifo.emptyB_0_cascade_\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__10042\,
            I => \N__10039\
        );

    \I__1391\ : InMux
    port map (
            O => \N__10039\,
            I => \N__10033\
        );

    \I__1390\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10033\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__10033\,
            I => \ufifo.tx_fsm.cstateZ0Z_1\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__10030\,
            I => \ufifo.tx_fsm.N_62_0_cascade_\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__10027\,
            I => \N__10020\
        );

    \I__1386\ : SRMux
    port map (
            O => \N__10026\,
            I => \N__10017\
        );

    \I__1385\ : CEMux
    port map (
            O => \N__10025\,
            I => \N__10014\
        );

    \I__1384\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10011\
        );

    \I__1383\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10008\
        );

    \I__1382\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10005\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__10017\,
            I => \N__10002\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__10014\,
            I => \N__9999\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__10011\,
            I => \N__9996\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__10008\,
            I => \N__9991\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10005\,
            I => \N__9991\
        );

    \I__1376\ : Span4Mux_h
    port map (
            O => \N__10002\,
            I => \N__9988\
        );

    \I__1375\ : Span4Mux_h
    port map (
            O => \N__9999\,
            I => \N__9985\
        );

    \I__1374\ : Span4Mux_h
    port map (
            O => \N__9996\,
            I => \N__9980\
        );

    \I__1373\ : Span4Mux_s2_v
    port map (
            O => \N__9991\,
            I => \N__9980\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__9988\,
            I => \ufifo.popFifo\
        );

    \I__1371\ : Odrv4
    port map (
            O => \N__9985\,
            I => \ufifo.popFifo\
        );

    \I__1370\ : Odrv4
    port map (
            O => \N__9980\,
            I => \ufifo.popFifo\
        );

    \I__1369\ : SRMux
    port map (
            O => \N__9973\,
            I => \N__9970\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__9970\,
            I => \N__9967\
        );

    \I__1367\ : Span4Mux_v
    port map (
            O => \N__9967\,
            I => \N__9963\
        );

    \I__1366\ : SRMux
    port map (
            O => \N__9966\,
            I => \N__9960\
        );

    \I__1365\ : Sp12to4
    port map (
            O => \N__9963\,
            I => \N__9956\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__9960\,
            I => \N__9953\
        );

    \I__1363\ : SRMux
    port map (
            O => \N__9959\,
            I => \N__9950\
        );

    \I__1362\ : Odrv12
    port map (
            O => \N__9956\,
            I => rst_i_3_i
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__9953\,
            I => rst_i_3_i
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__9950\,
            I => rst_i_3_i
        );

    \I__1359\ : InMux
    port map (
            O => \N__9943\,
            I => \N__9938\
        );

    \I__1358\ : InMux
    port map (
            O => \N__9942\,
            I => \N__9935\
        );

    \I__1357\ : InMux
    port map (
            O => \N__9941\,
            I => \N__9932\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__9938\,
            I => \N__9928\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__9935\,
            I => \N__9925\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__9932\,
            I => \N__9921\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__9931\,
            I => \N__9918\
        );

    \I__1352\ : Span4Mux_v
    port map (
            O => \N__9928\,
            I => \N__9911\
        );

    \I__1351\ : Span4Mux_v
    port map (
            O => \N__9925\,
            I => \N__9911\
        );

    \I__1350\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9908\
        );

    \I__1349\ : Span4Mux_v
    port map (
            O => \N__9921\,
            I => \N__9905\
        );

    \I__1348\ : InMux
    port map (
            O => \N__9918\,
            I => \N__9900\
        );

    \I__1347\ : InMux
    port map (
            O => \N__9917\,
            I => \N__9900\
        );

    \I__1346\ : InMux
    port map (
            O => \N__9916\,
            I => \N__9897\
        );

    \I__1345\ : Span4Mux_h
    port map (
            O => \N__9911\,
            I => \N__9892\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__9908\,
            I => \N__9892\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__9905\,
            I => \ufifo.emitcrlf_fsm.cstateZ0Z_0\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__9900\,
            I => \ufifo.emitcrlf_fsm.cstateZ0Z_0\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__9897\,
            I => \ufifo.emitcrlf_fsm.cstateZ0Z_0\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__9892\,
            I => \ufifo.emitcrlf_fsm.cstateZ0Z_0\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__9883\,
            I => \buart.Z_rx.bitcountlde_i_o2_0_cascade_\
        );

    \I__1338\ : InMux
    port map (
            O => \N__9880\,
            I => \N__9877\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__9877\,
            I => \N__9874\
        );

    \I__1336\ : Odrv12
    port map (
            O => \N__9874\,
            I => \Lab_UT.scdp.lsBitsi.q_esr_RNI0TMAZ0Z_3\
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__9871\,
            I => \Lab_UT.scdp.q_RNIRM8BD_3_cascade_\
        );

    \I__1334\ : InMux
    port map (
            O => \N__9868\,
            I => \N__9865\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__9865\,
            I => \N__9862\
        );

    \I__1332\ : Span4Mux_s3_h
    port map (
            O => \N__9862\,
            I => \N__9859\
        );

    \I__1331\ : Span4Mux_v
    port map (
            O => \N__9859\,
            I => \N__9856\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__9856\,
            I => \ufifo.txdataDZ0Z_3\
        );

    \I__1329\ : InMux
    port map (
            O => \N__9853\,
            I => \N__9850\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__9850\,
            I => \N__9845\
        );

    \I__1327\ : InMux
    port map (
            O => \N__9849\,
            I => \N__9842\
        );

    \I__1326\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9839\
        );

    \I__1325\ : Span12Mux_s10_v
    port map (
            O => \N__9845\,
            I => \N__9836\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__9842\,
            I => \N__9833\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__9839\,
            I => \Lab_UT.scdp.byteToDecrypt_0\
        );

    \I__1322\ : Odrv12
    port map (
            O => \N__9836\,
            I => \Lab_UT.scdp.byteToDecrypt_0\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__9833\,
            I => \Lab_UT.scdp.byteToDecrypt_0\
        );

    \I__1320\ : InMux
    port map (
            O => \N__9826\,
            I => \N__9821\
        );

    \I__1319\ : InMux
    port map (
            O => \N__9825\,
            I => \N__9818\
        );

    \I__1318\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9815\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__9821\,
            I => \Lab_UT.scdp.byteToDecrypt_3\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__9818\,
            I => \Lab_UT.scdp.byteToDecrypt_3\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__9815\,
            I => \Lab_UT.scdp.byteToDecrypt_3\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__9808\,
            I => \N__9805\
        );

    \I__1313\ : InMux
    port map (
            O => \N__9805\,
            I => \N__9802\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__9802\,
            I => \N__9799\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__9799\,
            I => \N__9794\
        );

    \I__1310\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9791\
        );

    \I__1309\ : InMux
    port map (
            O => \N__9797\,
            I => \N__9788\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__9794\,
            I => \ufifo.fifo.wraddrZ0Z_4\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__9791\,
            I => \ufifo.fifo.wraddrZ0Z_4\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__9788\,
            I => \ufifo.fifo.wraddrZ0Z_4\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__9781\,
            I => \N__9778\
        );

    \I__1304\ : InMux
    port map (
            O => \N__9778\,
            I => \N__9775\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__9775\,
            I => \N__9771\
        );

    \I__1302\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9767\
        );

    \I__1301\ : Span4Mux_v
    port map (
            O => \N__9771\,
            I => \N__9764\
        );

    \I__1300\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9761\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__9767\,
            I => \N__9758\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__9764\,
            I => \ufifo.fifo.rdaddrZ0Z_4\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__9761\,
            I => \ufifo.fifo.rdaddrZ0Z_4\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__9758\,
            I => \ufifo.fifo.rdaddrZ0Z_4\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__9751\,
            I => \N__9748\
        );

    \I__1294\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9745\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__9745\,
            I => \N__9741\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__9744\,
            I => \N__9737\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__9741\,
            I => \N__9734\
        );

    \I__1290\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9731\
        );

    \I__1289\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9728\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__9734\,
            I => \ufifo.fifo.wraddrZ0Z_5\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__9731\,
            I => \ufifo.fifo.wraddrZ0Z_5\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__9728\,
            I => \ufifo.fifo.wraddrZ0Z_5\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__9721\,
            I => \N__9718\
        );

    \I__1284\ : InMux
    port map (
            O => \N__9718\,
            I => \N__9715\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__9715\,
            I => \N__9711\
        );

    \I__1282\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9707\
        );

    \I__1281\ : Span12Mux_v
    port map (
            O => \N__9711\,
            I => \N__9704\
        );

    \I__1280\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9701\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__9707\,
            I => \N__9698\
        );

    \I__1278\ : Odrv12
    port map (
            O => \N__9704\,
            I => \ufifo.fifo.rdaddrZ0Z_5\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__9701\,
            I => \ufifo.fifo.rdaddrZ0Z_5\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__9698\,
            I => \ufifo.fifo.rdaddrZ0Z_5\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__9691\,
            I => \N__9688\
        );

    \I__1274\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9685\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__9685\,
            I => \N__9682\
        );

    \I__1272\ : Span4Mux_v
    port map (
            O => \N__9682\,
            I => \N__9677\
        );

    \I__1271\ : InMux
    port map (
            O => \N__9681\,
            I => \N__9674\
        );

    \I__1270\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9671\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__9677\,
            I => \ufifo.fifo.wraddrZ0Z_2\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__9674\,
            I => \ufifo.fifo.wraddrZ0Z_2\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__9671\,
            I => \ufifo.fifo.wraddrZ0Z_2\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__9664\,
            I => \N__9661\
        );

    \I__1265\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9658\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__9658\,
            I => \N__9654\
        );

    \I__1263\ : InMux
    port map (
            O => \N__9657\,
            I => \N__9650\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__9654\,
            I => \N__9647\
        );

    \I__1261\ : InMux
    port map (
            O => \N__9653\,
            I => \N__9644\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__9650\,
            I => \N__9641\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__9647\,
            I => \ufifo.fifo.rdaddrZ0Z_3\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__9644\,
            I => \ufifo.fifo.rdaddrZ0Z_3\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__9641\,
            I => \ufifo.fifo.rdaddrZ0Z_3\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__9634\,
            I => \N__9631\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9631\,
            I => \N__9628\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__9628\,
            I => \N__9624\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__9627\,
            I => \N__9620\
        );

    \I__1252\ : Span4Mux_v
    port map (
            O => \N__9624\,
            I => \N__9617\
        );

    \I__1251\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9614\
        );

    \I__1250\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9611\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__9617\,
            I => \ufifo.fifo.wraddrZ0Z_3\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__9614\,
            I => \ufifo.fifo.wraddrZ0Z_3\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__9611\,
            I => \ufifo.fifo.wraddrZ0Z_3\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__9604\,
            I => \N__9601\
        );

    \I__1245\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9598\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__9598\,
            I => \N__9594\
        );

    \I__1243\ : InMux
    port map (
            O => \N__9597\,
            I => \N__9590\
        );

    \I__1242\ : Span4Mux_v
    port map (
            O => \N__9594\,
            I => \N__9587\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9584\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__9590\,
            I => \N__9581\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__9587\,
            I => \ufifo.fifo.rdaddrZ0Z_2\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__9584\,
            I => \ufifo.fifo.rdaddrZ0Z_2\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__9581\,
            I => \ufifo.fifo.rdaddrZ0Z_2\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__9574\,
            I => \N__9571\
        );

    \I__1235\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9568\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__9568\,
            I => \N__9563\
        );

    \I__1233\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9560\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9557\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__9563\,
            I => \N__9550\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__9560\,
            I => \N__9550\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__9557\,
            I => \N__9550\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__9550\,
            I => \ufifo.fifo.wraddrZ0Z_1\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__9547\,
            I => \ufifo.fifo.un1_emptyB_NE_0_cascade_\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__9544\,
            I => \N__9541\
        );

    \I__1225\ : InMux
    port map (
            O => \N__9541\,
            I => \N__9538\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__9538\,
            I => \N__9534\
        );

    \I__1223\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9531\
        );

    \I__1222\ : Span4Mux_v
    port map (
            O => \N__9534\,
            I => \N__9527\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__9531\,
            I => \N__9524\
        );

    \I__1220\ : InMux
    port map (
            O => \N__9530\,
            I => \N__9521\
        );

    \I__1219\ : Span4Mux_v
    port map (
            O => \N__9527\,
            I => \N__9516\
        );

    \I__1218\ : Span4Mux_h
    port map (
            O => \N__9524\,
            I => \N__9516\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__9521\,
            I => \ufifo.fifo.rdaddrZ0Z_1\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__9516\,
            I => \ufifo.fifo.rdaddrZ0Z_1\
        );

    \I__1215\ : InMux
    port map (
            O => \N__9511\,
            I => \N__9507\
        );

    \I__1214\ : CascadeMux
    port map (
            O => \N__9510\,
            I => \N__9504\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__9507\,
            I => \N__9501\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9498\
        );

    \I__1211\ : Span4Mux_h
    port map (
            O => \N__9501\,
            I => \N__9495\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__9498\,
            I => \N__9492\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__9495\,
            I => \ufifo.tx_fsm.fifo_txdata_rdy\
        );

    \I__1208\ : Odrv12
    port map (
            O => \N__9492\,
            I => \ufifo.tx_fsm.fifo_txdata_rdy\
        );

    \I__1207\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9484\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__9484\,
            I => \N__9480\
        );

    \I__1205\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9477\
        );

    \I__1204\ : Odrv4
    port map (
            O => \N__9480\,
            I => \Lab_UT.scdp.e2dData_2\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__9477\,
            I => \Lab_UT.scdp.e2dData_2\
        );

    \I__1202\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9468\
        );

    \I__1201\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9465\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__9468\,
            I => \Lab_UT.scdp.N_59_i\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__9465\,
            I => \Lab_UT.scdp.N_59_i\
        );

    \I__1198\ : InMux
    port map (
            O => \N__9460\,
            I => \N__9457\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__9457\,
            I => \Lab_UT.scdp.pinst0.un12_pValidZ0Z_1\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9451\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__9451\,
            I => \N__9448\
        );

    \I__1194\ : Odrv12
    port map (
            O => \N__9448\,
            I => \Lab_UT.scdp.msBitsi.msBitsD_4\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9445\,
            I => \N__9439\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9444\,
            I => \N__9439\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__9439\,
            I => \N__9435\
        );

    \I__1190\ : InMux
    port map (
            O => \N__9438\,
            I => \N__9432\
        );

    \I__1189\ : Odrv12
    port map (
            O => \N__9435\,
            I => \Lab_UT.scdp.d2eData_3_4\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__9432\,
            I => \Lab_UT.scdp.d2eData_3_4\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__9427\,
            I => \Lab_UT.scdp.d2eData_3_4_cascade_\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__9424\,
            I => \Lab_UT.scdp.q_RNIIAV0D_0_cascade_\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9418\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__9418\,
            I => \Lab_UT.scdp.msBitsi.q_esr_RNI239EZ0Z_4\
        );

    \I__1183\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9412\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__9412\,
            I => \N__9409\
        );

    \I__1181\ : Span4Mux_v
    port map (
            O => \N__9409\,
            I => \N__9406\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__9406\,
            I => \ufifo.txdataDZ0Z_4\
        );

    \I__1179\ : InMux
    port map (
            O => \N__9403\,
            I => \N__9394\
        );

    \I__1178\ : InMux
    port map (
            O => \N__9402\,
            I => \N__9394\
        );

    \I__1177\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9394\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__9394\,
            I => \N__9390\
        );

    \I__1175\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9387\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__9390\,
            I => \Lab_UT.scdp.d2eData_3_3\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__9387\,
            I => \Lab_UT.scdp.d2eData_3_3\
        );

    \I__1172\ : InMux
    port map (
            O => \N__9382\,
            I => \N__9376\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9367\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9367\
        );

    \I__1169\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9367\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__9376\,
            I => \N__9364\
        );

    \I__1167\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9359\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9359\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__9367\,
            I => \N__9356\
        );

    \I__1164\ : Odrv12
    port map (
            O => \N__9364\,
            I => \Lab_UT.scdp.pValid_0\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__9359\,
            I => \Lab_UT.scdp.pValid_0\
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__9356\,
            I => \Lab_UT.scdp.pValid_0\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__9349\,
            I => \Lab_UT.scdp.d2eData_3_3_cascade_\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__9346\,
            I => \Lab_UT.scdp.d2eData_3_2_cascade_\
        );

    \I__1159\ : InMux
    port map (
            O => \N__9343\,
            I => \N__9340\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__9340\,
            I => \N__9337\
        );

    \I__1157\ : Span4Mux_h
    port map (
            O => \N__9337\,
            I => \N__9334\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__9334\,
            I => \Lab_UT.scdp.u2.byteToEncrypt_2\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__9331\,
            I => \N__9328\
        );

    \I__1154\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9319\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9327\,
            I => \N__9319\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9319\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__9319\,
            I => \Lab_UT.scdp.d2eData_2\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__9316\,
            I => \N__9312\
        );

    \I__1149\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9304\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9312\,
            I => \N__9304\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9304\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__9304\,
            I => \Lab_UT.scdp.d2eData_1\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__9301\,
            I => \N__9298\
        );

    \I__1144\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9295\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__9295\,
            I => \Lab_UT.scdp.lsBitsD_2\
        );

    \I__1142\ : InMux
    port map (
            O => \N__9292\,
            I => \N__9288\
        );

    \I__1141\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9285\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__9288\,
            I => \N__9282\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__9285\,
            I => \Lab_UT.scdp.d2eData_3_1\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__9282\,
            I => \Lab_UT.scdp.d2eData_3_1\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__9277\,
            I => \Lab_UT.scdp.pinst0.un12_pValidZ0Z_0_cascade_\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__9274\,
            I => \Lab_UT.scdp.un12_pValid_cascade_\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9267\
        );

    \I__1134\ : InMux
    port map (
            O => \N__9270\,
            I => \N__9264\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9267\,
            I => \N__9261\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__9264\,
            I => \N__9258\
        );

    \I__1131\ : Span12Mux_s11_v
    port map (
            O => \N__9261\,
            I => \N__9254\
        );

    \I__1130\ : Span4Mux_s3_h
    port map (
            O => \N__9258\,
            I => \N__9251\
        );

    \I__1129\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9248\
        );

    \I__1128\ : Odrv12
    port map (
            O => \N__9254\,
            I => \Lab_UT.scdp.d2eData_3_0\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__9251\,
            I => \Lab_UT.scdp.d2eData_3_0\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__9248\,
            I => \Lab_UT.scdp.d2eData_3_0\
        );

    \I__1125\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9238\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__9238\,
            I => \Lab_UT.scdp.un12_pValid\
        );

    \I__1123\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9229\
        );

    \I__1122\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9229\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__9229\,
            I => \N__9226\
        );

    \I__1120\ : Odrv12
    port map (
            O => \N__9226\,
            I => \Lab_UT.scdp.e2dData_6\
        );

    \I__1119\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9220\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__9220\,
            I => \N__9217\
        );

    \I__1117\ : Odrv12
    port map (
            O => \N__9217\,
            I => \Lab_UT.scdp.q_RNIDHFGA_3\
        );

    \I__1116\ : InMux
    port map (
            O => \N__9214\,
            I => \N__9211\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__9211\,
            I => \Lab_UT.scdp.d2eData_3_2\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9205\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__9205\,
            I => \N__9202\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__9202\,
            I => \N__9199\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__9199\,
            I => \Lab_UT.scdp.msBitsi.msBitsD_2\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__9196\,
            I => \Lab_UT.scdp.msBitsi.L4_tx_data_ns_1_2_cascade_\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9193\,
            I => \N__9190\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__9190\,
            I => \N__9187\
        );

    \I__1107\ : Span4Mux_s3_h
    port map (
            O => \N__9187\,
            I => \N__9184\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__9184\,
            I => \ufifo.txdataDZ0Z_2\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__9181\,
            I => \Lab_UT.scdp.d2eData_3_1_cascade_\
        );

    \I__1104\ : InMux
    port map (
            O => \N__9178\,
            I => \N__9175\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__9175\,
            I => \Lab_UT.scdp.q_RNIABC1D_1\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9172\,
            I => \N__9169\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__9169\,
            I => \N__9166\
        );

    \I__1100\ : Span4Mux_h
    port map (
            O => \N__9166\,
            I => \N__9163\
        );

    \I__1099\ : Odrv4
    port map (
            O => \N__9163\,
            I => \Lab_UT.scdp.u2.byteToEncrypt_1\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__9160\,
            I => \Lab_UT.scdp.d2eData_1_cascade_\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__9157\,
            I => \Lab_UT.scdp.lsBits_6_cascade_\
        );

    \I__1096\ : InMux
    port map (
            O => \N__9154\,
            I => \N__9151\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__9151\,
            I => \Lab_UT.scdp.lsBitsD_1\
        );

    \I__1094\ : InMux
    port map (
            O => \N__9148\,
            I => \N__9145\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__9145\,
            I => \N__9142\
        );

    \I__1092\ : Odrv12
    port map (
            O => \N__9142\,
            I => \Lab_UT.scdp.lsBitsi.lsBitsD_3\
        );

    \I__1091\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9130\
        );

    \I__1090\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9130\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9137\,
            I => \N__9130\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__9130\,
            I => \N__9127\
        );

    \I__1087\ : Span4Mux_h
    port map (
            O => \N__9127\,
            I => \N__9124\
        );

    \I__1086\ : Odrv4
    port map (
            O => \N__9124\,
            I => \Lab_UT.scdp.byteToEncrypt_3\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9118\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__9118\,
            I => \N__9115\
        );

    \I__1083\ : Span4Mux_v
    port map (
            O => \N__9115\,
            I => \N__9112\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__9112\,
            I => \Lab_UT.scdp.lsBitsD_6\
        );

    \I__1081\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9097\
        );

    \I__1080\ : InMux
    port map (
            O => \N__9108\,
            I => \N__9097\
        );

    \I__1079\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9097\
        );

    \I__1078\ : InMux
    port map (
            O => \N__9106\,
            I => \N__9097\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__9097\,
            I => \N__9094\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__9094\,
            I => \Lab_UT.scdp.d2eData_3_6\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__9091\,
            I => \Lab_UT.scdp.d2eData_3_6_cascade_\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9085\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9085\,
            I => \Lab_UT.scdp.u0.byteToDecrypt_6\
        );

    \I__1072\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9079\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__9079\,
            I => \N__9076\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__9076\,
            I => \N__9073\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__9073\,
            I => \ufifo.sb_ram512x8_inst_RNILSN11\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__9070\,
            I => \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0_cascade_\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9060\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9066\,
            I => \N__9060\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9065\,
            I => \N__9057\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__9060\,
            I => \N__9049\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__9049\
        );

    \I__1062\ : InMux
    port map (
            O => \N__9056\,
            I => \N__9044\
        );

    \I__1061\ : InMux
    port map (
            O => \N__9055\,
            I => \N__9041\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9054\,
            I => \N__9038\
        );

    \I__1059\ : Span4Mux_h
    port map (
            O => \N__9049\,
            I => \N__9035\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9048\,
            I => \N__9030\
        );

    \I__1057\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9030\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__9044\,
            I => ufifo_utb_txdata_sm0_0
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__9041\,
            I => ufifo_utb_txdata_sm0_0
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__9038\,
            I => ufifo_utb_txdata_sm0_0
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__9035\,
            I => ufifo_utb_txdata_sm0_0
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__9030\,
            I => ufifo_utb_txdata_sm0_0
        );

    \I__1051\ : InMux
    port map (
            O => \N__9019\,
            I => \N__9016\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__9016\,
            I => \N__9013\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__9013\,
            I => utb_txdata_2
        );

    \I__1048\ : InMux
    port map (
            O => \N__9010\,
            I => \N__9007\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__9007\,
            I => \N__9004\
        );

    \I__1046\ : Span12Mux_s3_h
    port map (
            O => \N__9004\,
            I => \N__9001\
        );

    \I__1045\ : Odrv12
    port map (
            O => \N__9001\,
            I => \ufifo.txdataDZ0Z_1\
        );

    \I__1044\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8995\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__8995\,
            I => \N__8992\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__8992\,
            I => \Lab_UT.scdp.msBitsi.msBitsD_1\
        );

    \I__1041\ : InMux
    port map (
            O => \N__8989\,
            I => \N__8986\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__8986\,
            I => \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8Z0Z_1\
        );

    \I__1039\ : InMux
    port map (
            O => \N__8983\,
            I => \N__8980\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__8980\,
            I => \N__8977\
        );

    \I__1037\ : Span4Mux_s3_h
    port map (
            O => \N__8977\,
            I => \N__8974\
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__8974\,
            I => \ufifo.txdataDZ0Z_5\
        );

    \I__1035\ : CEMux
    port map (
            O => \N__8971\,
            I => \N__8968\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__8968\,
            I => \N__8965\
        );

    \I__1033\ : Odrv12
    port map (
            O => \N__8965\,
            I => \Lab_UT.scdp.u2.sccEldByte_0\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__8962\,
            I => \Lab_UT.scdp.N_52_cascade_\
        );

    \I__1031\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8956\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__8956\,
            I => \Lab_UT.scdp.msBitsi.msBitsDZ0Z_0\
        );

    \I__1029\ : InMux
    port map (
            O => \N__8953\,
            I => \N__8947\
        );

    \I__1028\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8947\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__8947\,
            I => \N__8944\
        );

    \I__1026\ : Span4Mux_h
    port map (
            O => \N__8944\,
            I => \N__8941\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__8941\,
            I => \Lab_UT.scdp.byteToEncrypt_4\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__8938\,
            I => \N__8935\
        );

    \I__1023\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8932\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__8932\,
            I => \Lab_UT.scdp.b2a0.N_55\
        );

    \I__1021\ : InMux
    port map (
            O => \N__8929\,
            I => \N__8917\
        );

    \I__1020\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8917\
        );

    \I__1019\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8917\
        );

    \I__1018\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8917\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__8917\,
            I => \Lab_UT.scdp.d2eData_5\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__8914\,
            I => \Lab_UT.scdp.b2a0.N_55_cascade_\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__8911\,
            I => \Lab_UT.scdp.a2b.val_0_0Z0Z_3_cascade_\
        );

    \I__1014\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8905\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__8905\,
            I => \N__8902\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__8902\,
            I => \Lab_UT.scdp.msBitsi.q_esr_RNIF1M8Z0Z_6\
        );

    \I__1011\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8896\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__8896\,
            I => \Lab_UT.scdp.msBitsi.q_esr_RNIQQ8EZ0Z_0\
        );

    \I__1009\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8890\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__8890\,
            I => \N__8887\
        );

    \I__1007\ : Span4Mux_v
    port map (
            O => \N__8887\,
            I => \N__8884\
        );

    \I__1006\ : Odrv4
    port map (
            O => \N__8884\,
            I => \resetGen.escKey_0Z0Z_0\
        );

    \I__1005\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8878\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__8878\,
            I => \Lab_UT.scdp.msBitsi.msBitsD_6\
        );

    \I__1003\ : InMux
    port map (
            O => \N__8875\,
            I => \N__8872\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__8872\,
            I => \N__8869\
        );

    \I__1001\ : Span4Mux_v
    port map (
            O => \N__8869\,
            I => \N__8866\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__8866\,
            I => \Lab_UT.scdp.u2.byteToEncryptZ0Z_5\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__8863\,
            I => \Lab_UT.scdp.d2eData_5_cascade_\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__8860\,
            I => \N__8856\
        );

    \I__997\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8845\
        );

    \I__996\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8845\
        );

    \I__995\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8845\
        );

    \I__994\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8845\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__8845\,
            I => \N__8842\
        );

    \I__992\ : Span4Mux_v
    port map (
            O => \N__8842\,
            I => \N__8839\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__8839\,
            I => \Lab_UT.scdp.byteToEncrypt_6\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__8836\,
            I => \Lab_UT.scdp.q_RNI56C1D_0_cascade_\
        );

    \I__989\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8830\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__8830\,
            I => \ufifo.txdataDZ0Z_0\
        );

    \I__987\ : InMux
    port map (
            O => \N__8827\,
            I => \N__8824\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__8824\,
            I => \N__8821\
        );

    \I__985\ : Odrv4
    port map (
            O => \N__8821\,
            I => \ufifo.txdataDZ0Z_6\
        );

    \I__984\ : InMux
    port map (
            O => \N__8818\,
            I => \N__8813\
        );

    \I__983\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8808\
        );

    \I__982\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8808\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__8813\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__8808\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__8803\,
            I => \resetGen.reset_count_2_0_4_cascade_\
        );

    \I__978\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8797\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__8797\,
            I => \resetGen.un12_ci\
        );

    \I__976\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8791\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__8791\,
            I => \resetGen.un23_ci\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__8788\,
            I => \N__8785\
        );

    \I__973\ : InMux
    port map (
            O => \N__8785\,
            I => \N__8778\
        );

    \I__972\ : InMux
    port map (
            O => \N__8784\,
            I => \N__8773\
        );

    \I__971\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8773\
        );

    \I__970\ : InMux
    port map (
            O => \N__8782\,
            I => \N__8768\
        );

    \I__969\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8768\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__8778\,
            I => \N__8763\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__8773\,
            I => \N__8763\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__8768\,
            I => \N__8760\
        );

    \I__965\ : Span4Mux_h
    port map (
            O => \N__8763\,
            I => \N__8757\
        );

    \I__964\ : Span4Mux_h
    port map (
            O => \N__8760\,
            I => \N__8754\
        );

    \I__963\ : Odrv4
    port map (
            O => \N__8757\,
            I => \resetGen.escKeyZ0\
        );

    \I__962\ : Odrv4
    port map (
            O => \N__8754\,
            I => \resetGen.escKeyZ0\
        );

    \I__961\ : InMux
    port map (
            O => \N__8749\,
            I => \N__8743\
        );

    \I__960\ : InMux
    port map (
            O => \N__8748\,
            I => \N__8743\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__8743\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__958\ : InMux
    port map (
            O => \N__8740\,
            I => \bfn_4_4_0_\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__8737\,
            I => \resetGen.un12_ci_cascade_\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__8734\,
            I => \N__8731\
        );

    \I__955\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8728\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__8728\,
            I => \N__8724\
        );

    \I__953\ : InMux
    port map (
            O => \N__8727\,
            I => \N__8720\
        );

    \I__952\ : Span4Mux_v
    port map (
            O => \N__8724\,
            I => \N__8717\
        );

    \I__951\ : InMux
    port map (
            O => \N__8723\,
            I => \N__8714\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__8720\,
            I => \N__8711\
        );

    \I__949\ : Odrv4
    port map (
            O => \N__8717\,
            I => \ufifo.fifo.wraddrZ0Z_6\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__8714\,
            I => \ufifo.fifo.wraddrZ0Z_6\
        );

    \I__947\ : Odrv4
    port map (
            O => \N__8711\,
            I => \ufifo.fifo.wraddrZ0Z_6\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__8704\,
            I => \N__8701\
        );

    \I__945\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8698\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__8698\,
            I => \N__8694\
        );

    \I__943\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8690\
        );

    \I__942\ : Span4Mux_v
    port map (
            O => \N__8694\,
            I => \N__8687\
        );

    \I__941\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8684\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__8690\,
            I => \N__8681\
        );

    \I__939\ : Odrv4
    port map (
            O => \N__8687\,
            I => \ufifo.fifo.rdaddrZ0Z_7\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__8684\,
            I => \ufifo.fifo.rdaddrZ0Z_7\
        );

    \I__937\ : Odrv12
    port map (
            O => \N__8681\,
            I => \ufifo.fifo.rdaddrZ0Z_7\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__8674\,
            I => \N__8671\
        );

    \I__935\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8667\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__8670\,
            I => \N__8664\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__8667\,
            I => \N__8660\
        );

    \I__932\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8657\
        );

    \I__931\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8654\
        );

    \I__930\ : Span4Mux_v
    port map (
            O => \N__8660\,
            I => \N__8649\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__8657\,
            I => \N__8649\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__8654\,
            I => \ufifo.fifo.wraddrZ0Z_7\
        );

    \I__927\ : Odrv4
    port map (
            O => \N__8649\,
            I => \ufifo.fifo.wraddrZ0Z_7\
        );

    \I__926\ : CascadeMux
    port map (
            O => \N__8644\,
            I => \N__8641\
        );

    \I__925\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8638\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__8638\,
            I => \N__8635\
        );

    \I__923\ : Span4Mux_v
    port map (
            O => \N__8635\,
            I => \N__8630\
        );

    \I__922\ : InMux
    port map (
            O => \N__8634\,
            I => \N__8627\
        );

    \I__921\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8624\
        );

    \I__920\ : Sp12to4
    port map (
            O => \N__8630\,
            I => \N__8619\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__8627\,
            I => \N__8619\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__8624\,
            I => \ufifo.fifo.rdaddrZ0Z_6\
        );

    \I__917\ : Odrv12
    port map (
            O => \N__8619\,
            I => \ufifo.fifo.rdaddrZ0Z_6\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__8614\,
            I => \N__8611\
        );

    \I__915\ : InMux
    port map (
            O => \N__8611\,
            I => \N__8608\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__8608\,
            I => \N__8603\
        );

    \I__913\ : InMux
    port map (
            O => \N__8607\,
            I => \N__8600\
        );

    \I__912\ : InMux
    port map (
            O => \N__8606\,
            I => \N__8597\
        );

    \I__911\ : Span4Mux_v
    port map (
            O => \N__8603\,
            I => \N__8592\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__8600\,
            I => \N__8592\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__8597\,
            I => \ufifo.fifo.wraddrZ0Z_0\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__8592\,
            I => \ufifo.fifo.wraddrZ0Z_0\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__8587\,
            I => \N__8584\
        );

    \I__906\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8581\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__8581\,
            I => \N__8576\
        );

    \I__904\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8573\
        );

    \I__903\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8570\
        );

    \I__902\ : Sp12to4
    port map (
            O => \N__8576\,
            I => \N__8565\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__8573\,
            I => \N__8565\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8570\,
            I => \ufifo.fifo.rdaddrZ0Z_8\
        );

    \I__899\ : Odrv12
    port map (
            O => \N__8565\,
            I => \ufifo.fifo.rdaddrZ0Z_8\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__8560\,
            I => \N__8557\
        );

    \I__897\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8552\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__8556\,
            I => \N__8549\
        );

    \I__895\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8546\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__8552\,
            I => \N__8543\
        );

    \I__893\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8540\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__8546\,
            I => \N__8535\
        );

    \I__891\ : Span4Mux_v
    port map (
            O => \N__8543\,
            I => \N__8535\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__8540\,
            I => \N__8532\
        );

    \I__889\ : Odrv4
    port map (
            O => \N__8535\,
            I => \ufifo.fifo.wraddrZ0Z_8\
        );

    \I__888\ : Odrv4
    port map (
            O => \N__8532\,
            I => \ufifo.fifo.wraddrZ0Z_8\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__8527\,
            I => \N__8524\
        );

    \I__886\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8521\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__8521\,
            I => \N__8518\
        );

    \I__884\ : Span4Mux_v
    port map (
            O => \N__8518\,
            I => \N__8513\
        );

    \I__883\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8510\
        );

    \I__882\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8507\
        );

    \I__881\ : Sp12to4
    port map (
            O => \N__8513\,
            I => \N__8502\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__8510\,
            I => \N__8502\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__8507\,
            I => \ufifo.fifo.rdaddrZ0Z_0\
        );

    \I__878\ : Odrv12
    port map (
            O => \N__8502\,
            I => \ufifo.fifo.rdaddrZ0Z_0\
        );

    \I__877\ : InMux
    port map (
            O => \N__8497\,
            I => \N__8485\
        );

    \I__876\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8485\
        );

    \I__875\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8485\
        );

    \I__874\ : InMux
    port map (
            O => \N__8494\,
            I => \N__8485\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__8485\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__872\ : InMux
    port map (
            O => \N__8482\,
            I => \N__8473\
        );

    \I__871\ : InMux
    port map (
            O => \N__8481\,
            I => \N__8473\
        );

    \I__870\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8473\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__8473\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__868\ : InMux
    port map (
            O => \N__8470\,
            I => \bfn_4_2_0_\
        );

    \I__867\ : InMux
    port map (
            O => \N__8467\,
            I => \ufifo.fifo.un1_wraddr_cry_0\
        );

    \I__866\ : InMux
    port map (
            O => \N__8464\,
            I => \ufifo.fifo.un1_wraddr_cry_1\
        );

    \I__865\ : InMux
    port map (
            O => \N__8461\,
            I => \ufifo.fifo.un1_wraddr_cry_2\
        );

    \I__864\ : InMux
    port map (
            O => \N__8458\,
            I => \ufifo.fifo.un1_wraddr_cry_3\
        );

    \I__863\ : InMux
    port map (
            O => \N__8455\,
            I => \ufifo.fifo.un1_wraddr_cry_4\
        );

    \I__862\ : InMux
    port map (
            O => \N__8452\,
            I => \ufifo.fifo.un1_wraddr_cry_5\
        );

    \I__861\ : InMux
    port map (
            O => \N__8449\,
            I => \ufifo.fifo.un1_wraddr_cry_6\
        );

    \I__860\ : InMux
    port map (
            O => \N__8446\,
            I => \N__8443\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__8443\,
            I => \Lab_UT.scdp.u2.byteToEncrypt_0\
        );

    \I__858\ : InMux
    port map (
            O => \N__8440\,
            I => \ufifo.fifo.un1_rdaddr_cry_0\
        );

    \I__857\ : InMux
    port map (
            O => \N__8437\,
            I => \ufifo.fifo.un1_rdaddr_cry_1\
        );

    \I__856\ : InMux
    port map (
            O => \N__8434\,
            I => \ufifo.fifo.un1_rdaddr_cry_2\
        );

    \I__855\ : InMux
    port map (
            O => \N__8431\,
            I => \ufifo.fifo.un1_rdaddr_cry_3\
        );

    \I__854\ : InMux
    port map (
            O => \N__8428\,
            I => \ufifo.fifo.un1_rdaddr_cry_4\
        );

    \I__853\ : InMux
    port map (
            O => \N__8425\,
            I => \ufifo.fifo.un1_rdaddr_cry_5\
        );

    \I__852\ : InMux
    port map (
            O => \N__8422\,
            I => \ufifo.fifo.un1_rdaddr_cry_6\
        );

    \I__851\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8416\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__8416\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__849\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8410\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__8410\,
            I => \N__8407\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__8407\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__846\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8401\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__8401\,
            I => \N__8398\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__8398\,
            I => ufifo_utb_txdata_m0_4
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__8395\,
            I => \N__8392\
        );

    \I__842\ : InMux
    port map (
            O => \N__8392\,
            I => \N__8389\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__8389\,
            I => \N__8386\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__8386\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__839\ : CascadeMux
    port map (
            O => \N__8383\,
            I => \N__8380\
        );

    \I__838\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8377\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__8377\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__836\ : CEMux
    port map (
            O => \N__8374\,
            I => \N__8368\
        );

    \I__835\ : CEMux
    port map (
            O => \N__8373\,
            I => \N__8365\
        );

    \I__834\ : CEMux
    port map (
            O => \N__8372\,
            I => \N__8362\
        );

    \I__833\ : CEMux
    port map (
            O => \N__8371\,
            I => \N__8359\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__8368\,
            I => \N__8354\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8365\,
            I => \N__8354\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8362\,
            I => \N__8351\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__8359\,
            I => \N__8348\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__8354\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__827\ : Odrv4
    port map (
            O => \N__8351\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__8348\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__8341\,
            I => \N__8338\
        );

    \I__824\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8335\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__8335\,
            I => \N__8332\
        );

    \I__822\ : Odrv4
    port map (
            O => \N__8332\,
            I => \Lab_UT.scdp.byteToEncrypt_7\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__8329\,
            I => \ufifo.un4_rxDataValidNoEscZ0Z_1_cascade_\
        );

    \I__820\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8323\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__8323\,
            I => \ufifo.rxDataValidNoEscZ0\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__8320\,
            I => \N__8317\
        );

    \I__817\ : InMux
    port map (
            O => \N__8317\,
            I => \N__8314\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__8314\,
            I => \N__8311\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__8311\,
            I => \ufifo.fifo.fifo_txdata_3\
        );

    \I__814\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8305\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__8305\,
            I => \ufifo.fifo.fifo_txdata_4\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__8302\,
            I => \N__8299\
        );

    \I__811\ : InMux
    port map (
            O => \N__8299\,
            I => \N__8296\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__8296\,
            I => \N__8293\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__8293\,
            I => \ufifo.utb_txdata_m0_0\
        );

    \I__808\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__8287\,
            I => utb_txdata_0
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__8284\,
            I => \N__8281\
        );

    \I__805\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8275\
        );

    \I__804\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8275\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__8275\,
            I => \Lab_UT_dk_de_cr_2_reti\
        );

    \I__802\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8269\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__8269\,
            I => ufifo_utb_txdata_m0_3
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__8266\,
            I => \ufifo.sb_ram512x8_inst_RNIKRN11_cascade_\
        );

    \I__799\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8260\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__8260\,
            I => \ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0\
        );

    \I__797\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8254\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__8254\,
            I => utb_txdata_1
        );

    \I__795\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8248\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__8248\,
            I => \ufifo.fifo.fifo_txdata_0\
        );

    \I__793\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8242\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8239\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__8239\,
            I => \ufifo.fifo.fifo_txdata_6\
        );

    \I__790\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8233\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__8233\,
            I => \N__8230\
        );

    \I__788\ : Odrv4
    port map (
            O => \N__8230\,
            I => \ufifo.fifo.fifo_txdata_5\
        );

    \I__787\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8224\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__8224\,
            I => ufifo_utb_txdata_m0_5
        );

    \I__785\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8218\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__8218\,
            I => \ufifo.fifo.fifo_txdata_7\
        );

    \I__783\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8212\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__8212\,
            I => ufifo_utb_txdata_m0_7
        );

    \I__781\ : InMux
    port map (
            O => \N__8209\,
            I => \N__8206\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__8206\,
            I => ufifo_utb_txdata_m0_6
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__8203\,
            I => \N__8200\
        );

    \I__778\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8197\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__8197\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__8194\,
            I => \N__8191\
        );

    \I__775\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8188\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__8188\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__773\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8182\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8182\,
            I => \buart.Z_tx.counter_RNIVE1P1_1\
        );

    \I__771\ : InMux
    port map (
            O => \N__8179\,
            I => \buart.Z_tx.un1_bitcount_cry_0\
        );

    \I__770\ : InMux
    port map (
            O => \N__8176\,
            I => \N__8173\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__8173\,
            I => \buart.Z_tx.counter_RNIVE1P1_0_1\
        );

    \I__768\ : InMux
    port map (
            O => \N__8170\,
            I => \buart.Z_tx.un1_bitcount_cry_1\
        );

    \I__767\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__8164\,
            I => \buart.Z_tx.un1_bitcount_axb_3\
        );

    \I__765\ : InMux
    port map (
            O => \N__8161\,
            I => \buart.Z_tx.un1_bitcount_cry_2\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__8158\,
            I => \N__8155\
        );

    \I__763\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8152\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__8152\,
            I => \buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__8149\,
            I => \N__8146\
        );

    \I__760\ : InMux
    port map (
            O => \N__8146\,
            I => \N__8143\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__8143\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__758\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8135\
        );

    \I__757\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8130\
        );

    \I__756\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8130\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__8135\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__8130\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__753\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8122\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__8122\,
            I => \ufifo.fifo.fifo_txdata_2\
        );

    \I__751\ : InMux
    port map (
            O => \N__8119\,
            I => \N__8116\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__8116\,
            I => \ufifo.fifo.fifo_txdata_1\
        );

    \I__749\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8110\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__8110\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__747\ : IoInMux
    port map (
            O => \N__8107\,
            I => \N__8104\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__8104\,
            I => \N__8101\
        );

    \I__745\ : IoSpan4Mux
    port map (
            O => \N__8101\,
            I => \N__8098\
        );

    \I__744\ : Odrv4
    port map (
            O => \N__8098\,
            I => o_serial_data_c
        );

    \I__743\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8092\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__8092\,
            I => \uart_RXD\
        );

    \I__741\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8083\
        );

    \I__740\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8083\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__8083\,
            I => \N__8080\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__8080\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__737\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8074\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__8074\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__8071\,
            I => \N__8067\
        );

    \I__734\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8059\
        );

    \I__733\ : InMux
    port map (
            O => \N__8067\,
            I => \N__8059\
        );

    \I__732\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8059\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__8059\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__730\ : IoInMux
    port map (
            O => \N__8056\,
            I => \N__8053\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__8053\,
            I => \N__8050\
        );

    \I__728\ : IoSpan4Mux
    port map (
            O => \N__8050\,
            I => \N__8047\
        );

    \I__727\ : Span4Mux_s0_h
    port map (
            O => \N__8047\,
            I => \N__8044\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__8044\,
            I => \buart.Z_rx.N_41_i\
        );

    \I__725\ : InMux
    port map (
            O => \N__8041\,
            I => \N__8035\
        );

    \I__724\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8032\
        );

    \I__723\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8027\
        );

    \I__722\ : InMux
    port map (
            O => \N__8038\,
            I => \N__8027\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__8035\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__8032\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__8027\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__718\ : InMux
    port map (
            O => \N__8020\,
            I => \N__8017\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__8017\,
            I => \N__8014\
        );

    \I__716\ : Odrv4
    port map (
            O => \N__8014\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__8011\,
            I => \N__8006\
        );

    \I__714\ : InMux
    port map (
            O => \N__8010\,
            I => \N__8003\
        );

    \I__713\ : InMux
    port map (
            O => \N__8009\,
            I => \N__8000\
        );

    \I__712\ : InMux
    port map (
            O => \N__8006\,
            I => \N__7997\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__8003\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__8000\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__7997\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__708\ : InMux
    port map (
            O => \N__7990\,
            I => \N__7987\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__7987\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__706\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7981\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__7981\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__7978\,
            I => \N__7975\
        );

    \I__703\ : InMux
    port map (
            O => \N__7975\,
            I => \N__7970\
        );

    \I__702\ : InMux
    port map (
            O => \N__7974\,
            I => \N__7965\
        );

    \I__701\ : InMux
    port map (
            O => \N__7973\,
            I => \N__7965\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__7970\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__7965\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__698\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7954\
        );

    \I__697\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7947\
        );

    \I__696\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7947\
        );

    \I__695\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7947\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__7954\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__7947\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__7942\,
            I => \N__7938\
        );

    \I__691\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7935\
        );

    \I__690\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7932\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__7935\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__7932\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__687\ : InMux
    port map (
            O => \N__7927\,
            I => \N__7924\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__7924\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__685\ : InMux
    port map (
            O => \N__7921\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__684\ : InMux
    port map (
            O => \N__7918\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__683\ : InMux
    port map (
            O => \N__7915\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__682\ : InMux
    port map (
            O => \N__7912\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__681\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7903\
        );

    \I__680\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7903\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__7903\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__678\ : InMux
    port map (
            O => \N__7900\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__677\ : InMux
    port map (
            O => \N__7897\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__676\ : InMux
    port map (
            O => \N__7894\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__675\ : InMux
    port map (
            O => \N__7891\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__674\ : InMux
    port map (
            O => \N__7888\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__673\ : InMux
    port map (
            O => \N__7885\,
            I => \N__7879\
        );

    \I__672\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7879\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__7879\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__670\ : CascadeMux
    port map (
            O => \N__7876\,
            I => \N__7873\
        );

    \I__669\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7867\
        );

    \I__668\ : InMux
    port map (
            O => \N__7872\,
            I => \N__7867\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__7867\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__7864\,
            I => \N__7860\
        );

    \I__665\ : CascadeMux
    port map (
            O => \N__7863\,
            I => \N__7857\
        );

    \I__664\ : InMux
    port map (
            O => \N__7860\,
            I => \N__7852\
        );

    \I__663\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7852\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__7852\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__661\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7843\
        );

    \I__660\ : InMux
    port map (
            O => \N__7848\,
            I => \N__7843\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__7843\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__658\ : IoInMux
    port map (
            O => \N__7840\,
            I => \N__7837\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__7837\,
            I => \N__7834\
        );

    \I__656\ : Span12Mux_s1_v
    port map (
            O => \N__7834\,
            I => \N__7831\
        );

    \I__655\ : Span12Mux_v
    port map (
            O => \N__7831\,
            I => \N__7828\
        );

    \I__654\ : Odrv12
    port map (
            O => \N__7828\,
            I => \latticehx1k_pll_inst.clk\
        );

    \I__653\ : IoInMux
    port map (
            O => \N__7825\,
            I => \N__7822\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__7822\,
            I => \N__7819\
        );

    \I__651\ : IoSpan4Mux
    port map (
            O => \N__7819\,
            I => \N__7816\
        );

    \I__650\ : Odrv4
    port map (
            O => \N__7816\,
            I => clk_in_c
        );

    \IN_MUX_bfv_2_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_5_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_4_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_3_0_\
        );

    \IN_MUX_bfv_4_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ufifo.fifo.un1_wraddr_cry_7\,
            carryinitout => \bfn_4_4_0_\
        );

    \IN_MUX_bfv_4_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_1_0_\
        );

    \IN_MUX_bfv_4_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ufifo.fifo.un1_rdaddr_cry_7\,
            carryinitout => \bfn_4_2_0_\
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_4\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8056\,
            GLOBALBUFFEROUTPUT => \N_41_i_g\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7840\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12676\,
            GLOBALBUFFEROUTPUT => \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_g\
        );

    \resetGen.rst_0_iso_RNITVH4\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14086\,
            GLOBALBUFFEROUTPUT => \resetGen_rst_0_iso_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7960\,
            in2 => \N__7978\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7849\,
            in2 => \_gnd_net_\,
            in3 => \N__7900\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__22699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__12094\,
            in1 => \_gnd_net_\,
            in2 => \N__7876\,
            in3 => \N__7897\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__22699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7941\,
            in2 => \_gnd_net_\,
            in3 => \N__7894\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__22699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12095\,
            in1 => \N__7885\,
            in2 => \_gnd_net_\,
            in3 => \N__7891\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__22699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12093\,
            in2 => \N__7864\,
            in3 => \N__7888\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIGU38_6_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7884\,
            in1 => \N__7872\,
            in2 => \N__7863\,
            in3 => \N__7848\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__7959\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7974\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7958\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7973\,
            in1 => \N__7957\,
            in2 => \N__7942\,
            in3 => \N__7927\,
            lcout => \buart.Z_tx.N_255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1_0_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11374\,
            in1 => \N__9917\,
            in2 => \_gnd_net_\,
            in3 => \N__11462\,
            lcout => \ufifo.crlfdone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_0_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__11463\,
            in1 => \N__11375\,
            in2 => \N__9931\,
            in3 => \N__20243\,
            lcout => \ufifo.emitcrlf_fsm.cstateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8039\,
            in2 => \N__8071\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8139\,
            in2 => \_gnd_net_\,
            in3 => \N__7921\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10367\,
            in1 => \N__7909\,
            in2 => \_gnd_net_\,
            in3 => \N__7918\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__22689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8009\,
            in2 => \_gnd_net_\,
            in3 => \N__7915\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__8089\,
            in1 => \N__10366\,
            in2 => \N__10182\,
            in3 => \N__7912\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7908\,
            in1 => \N__8138\,
            in2 => \N__8011\,
            in3 => \N__8066\,
            lcout => \buart.Z_rx.Z_baudgen.ser_clk_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8088\,
            in1 => \N__8038\,
            in2 => \_gnd_net_\,
            in3 => \N__8077\,
            lcout => \buart.Z_rx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10365\,
            in1 => \N__8041\,
            in2 => \_gnd_net_\,
            in3 => \N__8070\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_4_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__10170\,
            in1 => \N__10497\,
            in2 => \N__10408\,
            in3 => \N__10609\,
            lcout => \buart.Z_rx.N_41_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8040\,
            in2 => \_gnd_net_\,
            in3 => \N__10377\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__10171\,
            in1 => \N__8020\,
            in2 => \N__10378\,
            in3 => \N__8010\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_0_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111111111"
        )
    port map (
            in0 => \N__11386\,
            in1 => \N__9924\,
            in2 => \_gnd_net_\,
            in3 => \N__11467\,
            lcout => ufifo_utb_txdata_sm0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7990\,
            in1 => \N__8290\,
            in2 => \_gnd_net_\,
            in3 => \N__12038\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22676\,
            ce => \N__8374\,
            sr => \N__18063\
        );

    \buart.Z_tx.shifter_6_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__8227\,
            in1 => \N__9055\,
            in2 => \N__8194\,
            in3 => \N__12039\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22676\,
            ce => \N__8374\,
            sr => \N__18063\
        );

    \buart.Z_tx.shifter_2_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12037\,
            in1 => \N__8413\,
            in2 => \_gnd_net_\,
            in3 => \N__8257\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22676\,
            ce => \N__8374\,
            sr => \N__18063\
        );

    \buart.Z_tx.shifter_0_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7984\,
            in2 => \_gnd_net_\,
            in3 => \N__12051\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22668\,
            ce => \N__8371\,
            sr => \N__18065\
        );

    \buart.Z_tx.uart_tx_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__12050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8113\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22668\,
            ce => \N__8371\,
            sr => \N__18065\
        );

    \buart.Z_rx.hh_1_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10212\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22664\,
            ce => 'H',
            sr => \N__18066\
        );

    \buart.Z_rx.hh_0_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8095\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22655\,
            ce => 'H',
            sr => \N__18067\
        );

    \ufifo.tx_fsm.cstate_3_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10024\,
            lcout => \ufifo.tx_fsm.fifo_txdata_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22697\,
            ce => 'H',
            sr => \N__9959\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_1_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12086\,
            in2 => \_gnd_net_\,
            in3 => \N__12176\,
            lcout => \buart.Z_tx.counter_RNIVE1P1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_0_1_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__12177\,
            in1 => \_gnd_net_\,
            in2 => \N__12103\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.counter_RNIVE1P1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.state_ret_5_RNIAFUE_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20271\,
            lcout => rst_i_3_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__12178\,
            in1 => \_gnd_net_\,
            in2 => \N__12104\,
            in3 => \N__10095\,
            lcout => \buart.Z_tx.un1_bitcount_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.un1_bitcount_cry_0_0_c_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11968\,
            in2 => \N__8158\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_5_0_\,
            carryout => \buart.Z_tx.un1_bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_1_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__12048\,
            in1 => \N__8185\,
            in2 => \N__10117\,
            in3 => \N__8179\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \buart.Z_tx.un1_bitcount_cry_0\,
            carryout => \buart.Z_tx.un1_bitcount_cry_1\,
            clk => \N__22690\,
            ce => 'H',
            sr => \N__18070\
        );

    \buart.Z_tx.bitcount_2_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__12047\,
            in1 => \N__8176\,
            in2 => \N__10135\,
            in3 => \N__8170\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.un1_bitcount_cry_1\,
            carryout => \buart.Z_tx.un1_bitcount_cry_2\,
            clk => \N__22690\,
            ce => 'H',
            sr => \N__18070\
        );

    \buart.Z_tx.bitcount_3_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__12049\,
            in1 => \N__8167\,
            in2 => \_gnd_net_\,
            in3 => \N__8161\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22690\,
            ce => 'H',
            sr => \N__18070\
        );

    \resetGen.rst_0_iso_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22761\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \resetGen_rst_0_iso\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.un1_bitcount_cry_0_0_c_RNO_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12096\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12158\,
            lcout => \buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__10364\,
            in1 => \N__8140\,
            in2 => \N__8149\,
            in3 => \N__10178\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__11387\,
            in1 => \N__9916\,
            in2 => \_gnd_net_\,
            in3 => \N__11469\,
            lcout => \ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNILSN11_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11242\,
            in1 => \N__8125\,
            in2 => \_gnd_net_\,
            in3 => \N__15686\,
            lcout => \ufifo.sb_ram512x8_inst_RNILSN11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNIKRN11_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15771\,
            in1 => \N__11262\,
            in2 => \_gnd_net_\,
            in3 => \N__8119\,
            lcout => OPEN,
            ltout => \ufifo.sb_ram512x8_inst_RNIKRN11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIQ6FP3_0_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__9048\,
            in1 => \_gnd_net_\,
            in2 => \N__8266\,
            in3 => \N__8263\,
            lcout => utb_txdata_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNIJQN11_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11263\,
            in1 => \N__8251\,
            in2 => \_gnd_net_\,
            in3 => \N__16166\,
            lcout => \ufifo.utb_txdata_m0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNIP0O11_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8245\,
            in1 => \N__11267\,
            in2 => \_gnd_net_\,
            in3 => \N__17074\,
            lcout => ufifo_utb_txdata_m0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNIA4BA7_3_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001100"
        )
    port map (
            in0 => \N__11264\,
            in1 => \N__9047\,
            in2 => \N__9510\,
            in3 => \N__8326\,
            lcout => ufifo_utb_txdata_rdy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNIOVN11_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8236\,
            in1 => \N__11266\,
            in2 => \_gnd_net_\,
            in3 => \N__13437\,
            lcout => ufifo_utb_txdata_m0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNIQ1O11_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8221\,
            in1 => \N__11265\,
            in2 => \_gnd_net_\,
            in3 => \N__16964\,
            lcout => ufifo_utb_txdata_m0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_8_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__8215\,
            in1 => \N__9054\,
            in2 => \_gnd_net_\,
            in3 => \N__12036\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22669\,
            ce => \N__8373\,
            sr => \N__18064\
        );

    \buart.Z_tx.shifter_7_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__12035\,
            in1 => \N__8209\,
            in2 => \N__8203\,
            in3 => \N__9056\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22669\,
            ce => \N__8373\,
            sr => \N__18064\
        );

    \ufifo.un4_rxDataValidNoEsc_1_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__13318\,
            in1 => \N__16955\,
            in2 => \N__15702\,
            in3 => \N__11680\,
            lcout => OPEN,
            ltout => \ufifo.un4_rxDataValidNoEscZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.rxDataValidNoEsc_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100000000"
        )
    port map (
            in0 => \N__11592\,
            in1 => \N__8280\,
            in2 => \N__8329\,
            in3 => \N__20809\,
            lcout => \ufifo.rxDataValidNoEscZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__20810\,
            in1 => \N__8893\,
            in2 => \N__8284\,
            in3 => \N__11593\,
            lcout => \resetGen.escKeyZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_3_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11041\,
            in1 => \N__10798\,
            in2 => \N__8341\,
            in3 => \N__10954\,
            lcout => \Lab_UT.scdp.N_48_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNIMTN11_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__11922\,
            in1 => \_gnd_net_\,
            in2 => \N__8320\,
            in3 => \N__11268\,
            lcout => ufifo_utb_txdata_m0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.sb_ram512x8_inst_RNINUN11_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11269\,
            in1 => \N__8308\,
            in2 => \_gnd_net_\,
            in3 => \N__13377\,
            lcout => ufifo_utb_txdata_m0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNI6GJD2_0_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110000"
        )
    port map (
            in0 => \N__11394\,
            in1 => \N__9941\,
            in2 => \N__8302\,
            in3 => \N__11473\,
            lcout => utb_txdata_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_2_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11921\,
            in2 => \_gnd_net_\,
            in3 => \N__13376\,
            lcout => \Lab_UT_dk_de_cr_2_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI9JC39_1_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__12179\,
            in1 => \N__12105\,
            in2 => \_gnd_net_\,
            in3 => \N__12040\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_4_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010111011"
        )
    port map (
            in0 => \N__8272\,
            in1 => \N__9066\,
            in2 => \N__8383\,
            in3 => \N__12042\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22656\,
            ce => \N__8372\,
            sr => \N__18068\
        );

    \buart.Z_tx.shifter_3_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12041\,
            in1 => \N__8419\,
            in2 => \_gnd_net_\,
            in3 => \N__9019\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22656\,
            ce => \N__8372\,
            sr => \N__18068\
        );

    \buart.Z_tx.shifter_5_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__8404\,
            in1 => \N__9067\,
            in2 => \N__8395\,
            in3 => \N__12043\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22656\,
            ce => \N__8372\,
            sr => \N__18068\
        );

    \Lab_UT.scdp.u2.q_esr_1_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15782\,
            lcout => \Lab_UT.scdp.u2.byteToEncrypt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22651\,
            ce => \N__8971\,
            sr => \N__18039\
        );

    \Lab_UT.scdp.u2.q_esr_2_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15687\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scdp.u2.byteToEncrypt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22651\,
            ce => \N__8971\,
            sr => \N__18039\
        );

    \Lab_UT.scdp.u2.q_esr_3_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11934\,
            lcout => \Lab_UT.scdp.byteToEncrypt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22651\,
            ce => \N__8971\,
            sr => \N__18039\
        );

    \Lab_UT.scdp.u2.q_esr_4_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13378\,
            lcout => \Lab_UT.scdp.byteToEncrypt_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22651\,
            ce => \N__8971\,
            sr => \N__18039\
        );

    \Lab_UT.scdp.u2.q_esr_5_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13438\,
            lcout => \Lab_UT.scdp.u2.byteToEncryptZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22651\,
            ce => \N__8971\,
            sr => \N__18039\
        );

    \Lab_UT.scdp.u2.q_esr_6_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17075\,
            lcout => \Lab_UT.scdp.byteToEncrypt_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22651\,
            ce => \N__8971\,
            sr => \N__18039\
        );

    \Lab_UT.scdp.u2.q_esr_7_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16965\,
            lcout => \Lab_UT.scdp.byteToEncrypt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22651\,
            ce => \N__8971\,
            sr => \N__18039\
        );

    \Lab_UT.scdp.u2.q_esr_0_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16167\,
            lcout => \Lab_UT.scdp.u2.byteToEncrypt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22651\,
            ce => \N__8971\,
            sr => \N__18039\
        );

    \Lab_UT.scdp.u2.q_esr_RNIT8JT_0_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8446\,
            in2 => \_gnd_net_\,
            in3 => \N__9270\,
            lcout => \Lab_UT.scdp.d2eData_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.rdaddr_0_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8516\,
            in2 => \N__10027\,
            in3 => \N__10023\,
            lcout => \ufifo.fifo.rdaddrZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_1_0_\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_0\,
            clk => \N__22698\,
            ce => 'H',
            sr => \N__18050\
        );

    \ufifo.fifo.rdaddr_1_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9530\,
            in2 => \_gnd_net_\,
            in3 => \N__8440\,
            lcout => \ufifo.fifo.rdaddrZ0Z_1\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_0\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_1\,
            clk => \N__22698\,
            ce => 'H',
            sr => \N__18050\
        );

    \ufifo.fifo.rdaddr_2_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9593\,
            in2 => \_gnd_net_\,
            in3 => \N__8437\,
            lcout => \ufifo.fifo.rdaddrZ0Z_2\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_1\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_2\,
            clk => \N__22698\,
            ce => 'H',
            sr => \N__18050\
        );

    \ufifo.fifo.rdaddr_3_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9653\,
            in2 => \_gnd_net_\,
            in3 => \N__8434\,
            lcout => \ufifo.fifo.rdaddrZ0Z_3\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_2\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_3\,
            clk => \N__22698\,
            ce => 'H',
            sr => \N__18050\
        );

    \ufifo.fifo.rdaddr_4_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9770\,
            in2 => \_gnd_net_\,
            in3 => \N__8431\,
            lcout => \ufifo.fifo.rdaddrZ0Z_4\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_3\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_4\,
            clk => \N__22698\,
            ce => 'H',
            sr => \N__18050\
        );

    \ufifo.fifo.rdaddr_5_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9710\,
            in2 => \_gnd_net_\,
            in3 => \N__8428\,
            lcout => \ufifo.fifo.rdaddrZ0Z_5\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_4\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_5\,
            clk => \N__22698\,
            ce => 'H',
            sr => \N__18050\
        );

    \ufifo.fifo.rdaddr_6_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8633\,
            in2 => \_gnd_net_\,
            in3 => \N__8425\,
            lcout => \ufifo.fifo.rdaddrZ0Z_6\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_5\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_6\,
            clk => \N__22698\,
            ce => 'H',
            sr => \N__18050\
        );

    \ufifo.fifo.rdaddr_7_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8693\,
            in2 => \_gnd_net_\,
            in3 => \N__8422\,
            lcout => \ufifo.fifo.rdaddrZ0Z_7\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_rdaddr_cry_6\,
            carryout => \ufifo.fifo.un1_rdaddr_cry_7\,
            clk => \N__22698\,
            ce => 'H',
            sr => \N__18050\
        );

    \ufifo.fifo.rdaddr_8_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8579\,
            in2 => \_gnd_net_\,
            in3 => \N__8470\,
            lcout => \ufifo.fifo.rdaddrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22694\,
            ce => 'H',
            sr => \N__18047\
        );

    \ufifo.fifo.wraddr_0_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8606\,
            in2 => \N__11090\,
            in3 => \N__11083\,
            lcout => \ufifo.fifo.wraddrZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_3_0_\,
            carryout => \ufifo.fifo.un1_wraddr_cry_0\,
            clk => \N__22691\,
            ce => 'H',
            sr => \N__18045\
        );

    \ufifo.fifo.wraddr_1_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9567\,
            in2 => \_gnd_net_\,
            in3 => \N__8467\,
            lcout => \ufifo.fifo.wraddrZ0Z_1\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_0\,
            carryout => \ufifo.fifo.un1_wraddr_cry_1\,
            clk => \N__22691\,
            ce => 'H',
            sr => \N__18045\
        );

    \ufifo.fifo.wraddr_2_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9681\,
            in2 => \_gnd_net_\,
            in3 => \N__8464\,
            lcout => \ufifo.fifo.wraddrZ0Z_2\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_1\,
            carryout => \ufifo.fifo.un1_wraddr_cry_2\,
            clk => \N__22691\,
            ce => 'H',
            sr => \N__18045\
        );

    \ufifo.fifo.wraddr_3_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9623\,
            in2 => \_gnd_net_\,
            in3 => \N__8461\,
            lcout => \ufifo.fifo.wraddrZ0Z_3\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_2\,
            carryout => \ufifo.fifo.un1_wraddr_cry_3\,
            clk => \N__22691\,
            ce => 'H',
            sr => \N__18045\
        );

    \ufifo.fifo.wraddr_4_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9798\,
            in2 => \_gnd_net_\,
            in3 => \N__8458\,
            lcout => \ufifo.fifo.wraddrZ0Z_4\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_3\,
            carryout => \ufifo.fifo.un1_wraddr_cry_4\,
            clk => \N__22691\,
            ce => 'H',
            sr => \N__18045\
        );

    \ufifo.fifo.wraddr_5_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9740\,
            in2 => \_gnd_net_\,
            in3 => \N__8455\,
            lcout => \ufifo.fifo.wraddrZ0Z_5\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_4\,
            carryout => \ufifo.fifo.un1_wraddr_cry_5\,
            clk => \N__22691\,
            ce => 'H',
            sr => \N__18045\
        );

    \ufifo.fifo.wraddr_6_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8723\,
            in2 => \_gnd_net_\,
            in3 => \N__8452\,
            lcout => \ufifo.fifo.wraddrZ0Z_6\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_5\,
            carryout => \ufifo.fifo.un1_wraddr_cry_6\,
            clk => \N__22691\,
            ce => 'H',
            sr => \N__18045\
        );

    \ufifo.fifo.wraddr_7_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8663\,
            in2 => \_gnd_net_\,
            in3 => \N__8449\,
            lcout => \ufifo.fifo.wraddrZ0Z_7\,
            ltout => OPEN,
            carryin => \ufifo.fifo.un1_wraddr_cry_6\,
            carryout => \ufifo.fifo.un1_wraddr_cry_7\,
            clk => \N__22691\,
            ce => 'H',
            sr => \N__18045\
        );

    \ufifo.fifo.wraddr_8_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8555\,
            in2 => \_gnd_net_\,
            in3 => \N__8740\,
            lcout => \ufifo.fifo.wraddrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22684\,
            ce => 'H',
            sr => \N__18043\
        );

    \resetGen.uu0.counter_gen_label_3__un23_ci_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8480\,
            in1 => \N__8495\,
            in2 => \_gnd_net_\,
            in3 => \N__8816\,
            lcout => \resetGen.un23_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__8496\,
            in1 => \N__22764\,
            in2 => \_gnd_net_\,
            in3 => \N__8783\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22677\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_2__un12_ci_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8481\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8494\,
            lcout => \resetGen.un12_ci\,
            ltout => \resetGen.un12_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011010"
        )
    port map (
            in0 => \N__8817\,
            in1 => \N__22763\,
            in2 => \N__8737\,
            in3 => \N__8784\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22677\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_RNI8A8U_6_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__8727\,
            in1 => \N__8697\,
            in2 => \N__8670\,
            in3 => \N__8634\,
            lcout => \ufifo.fifo.un1_emptyB_NE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_RNIUV7U_8_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__8607\,
            in1 => \N__8580\,
            in2 => \N__8556\,
            in3 => \N__8517\,
            lcout => \ufifo.fifo.un1_emptyB_NE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_10_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011111"
        )
    port map (
            in0 => \N__18441\,
            in1 => \N__18946\,
            in2 => \N__17615\,
            in3 => \N__20098\,
            lcout => \Lab_UT.scctrl.g0_7_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000110"
        )
    port map (
            in0 => \N__8497\,
            in1 => \N__8482\,
            in2 => \N__8788\,
            in3 => \N__22765\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22677\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNI56C1D_0_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__9853\,
            in1 => \N__9271\,
            in2 => \_gnd_net_\,
            in3 => \N__9382\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.q_RNI56C1D_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_0_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8899\,
            in2 => \N__8836\,
            in3 => \N__17838\,
            lcout => \ufifo.txdataDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIQOQA1_0_3_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11432\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart__tx_uart_busy_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_6_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8908\,
            in1 => \N__17839\,
            in2 => \_gnd_net_\,
            in3 => \N__9223\,
            lcout => \ufifo.txdataDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNO_0_4_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8748\,
            in2 => \_gnd_net_\,
            in3 => \N__8818\,
            lcout => OPEN,
            ltout => \resetGen.reset_count_2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__8781\,
            in1 => \N__22744\,
            in2 => \N__8803\,
            in3 => \N__8800\,
            lcout => rst_i_3_reti,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000110"
        )
    port map (
            in0 => \N__8794\,
            in1 => \N__8749\,
            in2 => \N__22766\,
            in3 => \N__8782\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_3_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__21546\,
            in1 => \N__21489\,
            in2 => \N__20272\,
            in3 => \N__14545\,
            lcout => \Lab_UT.scctrl.next_state_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22665\,
            ce => \N__14793\,
            sr => \N__18071\
        );

    \Lab_UT.scdp.lsBitsi.q_esr_RNI0TMA_3_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9148\,
            in1 => \N__12208\,
            in2 => \_gnd_net_\,
            in3 => \N__18164\,
            lcout => \Lab_UT.scdp.lsBitsi.q_esr_RNI0TMAZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNIF1M8_6_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18165\,
            in1 => \N__8881\,
            in2 => \_gnd_net_\,
            in3 => \N__9121\,
            lcout => \Lab_UT.scdp.msBitsi.q_esr_RNIF1M8Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNIQQ8E_0_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8959\,
            in1 => \N__12337\,
            in2 => \_gnd_net_\,
            in3 => \N__18166\,
            lcout => \Lab_UT.scdp.msBitsi.q_esr_RNIQQ8EZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIOP0V3_4_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10197\,
            in2 => \_gnd_net_\,
            in3 => \N__20808\,
            lcout => \buart.Z_rx.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_0_0_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__16774\,
            in1 => \N__15695\,
            in2 => \_gnd_net_\,
            in3 => \N__16943\,
            lcout => \resetGen.escKey_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_2_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001011001000"
        )
    port map (
            in0 => \N__8927\,
            in1 => \N__9109\,
            in2 => \N__8938\,
            in3 => \N__8855\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22657\,
            ce => \N__13200\,
            sr => \N__18038\
        );

    \Lab_UT.scdp.msBitsi.q_esr_6_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100010010"
        )
    port map (
            in0 => \N__9107\,
            in1 => \N__12259\,
            in2 => \N__8860\,
            in3 => \N__8928\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22657\,
            ce => \N__13200\,
            sr => \N__18038\
        );

    \Lab_UT.scdp.msBitsi.q_esr_4_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110001"
        )
    port map (
            in0 => \N__8929\,
            in1 => \N__9108\,
            in2 => \N__12267\,
            in3 => \N__8859\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22657\,
            ce => \N__13200\,
            sr => \N__18038\
        );

    \Lab_UT.scdp.u2.q_esr_RNIKRG71_5_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8875\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10852\,
            lcout => \Lab_UT.scdp.d2eData_5\,
            ltout => \Lab_UT.scdp.d2eData_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.b2a0.asciiHex_2_i_o3_3_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9106\,
            in2 => \N__8863\,
            in3 => \N__8854\,
            lcout => \Lab_UT.scdp.N_52\,
            ltout => \Lab_UT.scdp.N_52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_0_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010010110"
        )
    port map (
            in0 => \N__9445\,
            in1 => \N__8953\,
            in2 => \N__8962\,
            in3 => \N__12263\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22657\,
            ce => \N__13200\,
            sr => \N__18038\
        );

    \Lab_UT.scdp.b2a0.asciiHex_2_0_a2_0_o2_0_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111101110"
        )
    port map (
            in0 => \N__8952\,
            in1 => \N__12258\,
            in2 => \_gnd_net_\,
            in3 => \N__9444\,
            lcout => \Lab_UT.scdp.b2a0.N_55\,
            ltout => \Lab_UT.scdp.b2a0.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_1_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8926\,
            in2 => \N__8914\,
            in3 => \N__12219\,
            lcout => \Lab_UT.scdp.msBitsi.msBitsD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22657\,
            ce => \N__13200\,
            sr => \N__18038\
        );

    \Lab_UT.scctrl.g0_17_N_2L1_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10599\,
            in1 => \N__12424\,
            in2 => \N__16505\,
            in3 => \N__10650\,
            lcout => \Lab_UT.scctrl.g0_17_N_2LZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_fast_RNI1CIH1_2_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__12423\,
            in1 => \N__10649\,
            in2 => \N__16504\,
            in3 => \N__10598\,
            lcout => \buart.Z_rx.shifter_0_fast_RNI1CIH1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_fast_2_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11925\,
            lcout => \buart__rx_shifter_0_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22652\,
            ce => \N__16752\,
            sr => \N__18072\
        );

    \buart.Z_rx.shifter_ret_1_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15694\,
            lcout => bu_rx_data_i_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22652\,
            ce => \N__16752\,
            sr => \N__18072\
        );

    \Lab_UT.scdp.a2b.val_0_0_3_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000000"
        )
    port map (
            in0 => \N__11923\,
            in1 => \N__16169\,
            in2 => \N__15704\,
            in3 => \N__14845\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.a2b.val_0_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.val_0_3_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11626\,
            in2 => \N__8911\,
            in3 => \N__11924\,
            lcout => \Lab_UT.scdp.val_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.val18_1_i_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16168\,
            in2 => \_gnd_net_\,
            in3 => \N__14844\,
            lcout => \N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIM7051_14_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10840\,
            in1 => \N__10677\,
            in2 => \N__11797\,
            in3 => \N__11824\,
            lcout => \Lab_UT.scdp.d2eData_3_6\,
            ltout => \Lab_UT.scdp.d2eData_3_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_esr_RNIA29D1_2_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9091\,
            in3 => \N__9088\,
            lcout => \Lab_UT.scdp.e2dData_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_esr_2_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__15696\,
            in1 => \N__15772\,
            in2 => \_gnd_net_\,
            in3 => \N__15818\,
            lcout => \Lab_UT.scdp.u0.byteToDecrypt_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22645\,
            ce => \N__13126\,
            sr => \N__18040\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2_0_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11395\,
            in1 => \N__9942\,
            in2 => \_gnd_net_\,
            in3 => \N__11468\,
            lcout => OPEN,
            ltout => \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNIR7FP3_0_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9082\,
            in2 => \N__9070\,
            in3 => \N__9065\,
            lcout => utb_txdata_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_1_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8989\,
            in1 => \N__17830\,
            in2 => \_gnd_net_\,
            in3 => \N__9178\,
            lcout => \ufifo.txdataDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8_1_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8998\,
            in1 => \N__9154\,
            in2 => \_gnd_net_\,
            in3 => \N__18155\,
            lcout => \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_5_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__9381\,
            in1 => \N__17832\,
            in2 => \N__13156\,
            in3 => \N__11191\,
            lcout => \ufifo.txdataDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u2.q_esr_ctle_7_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18091\,
            in2 => \_gnd_net_\,
            in3 => \N__12823\,
            lcout => \Lab_UT.scdp.u2.sccEldByte_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNI7PL8_2_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__18156\,
            in1 => \_gnd_net_\,
            in2 => \N__9301\,
            in3 => \N__9208\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.msBitsi.L4_tx_data_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_2_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101001001110"
        )
    port map (
            in0 => \N__17831\,
            in1 => \N__9487\,
            in2 => \N__9196\,
            in3 => \N__9380\,
            lcout => \ufifo.txdataDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNID22R_1_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10737\,
            in1 => \N__10689\,
            in2 => \N__10813\,
            in3 => \N__12526\,
            lcout => \Lab_UT.scdp.d2eData_3_1\,
            ltout => \Lab_UT.scdp.d2eData_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNIABC1D_1_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14002\,
            in2 => \N__9181\,
            in3 => \N__9379\,
            lcout => \Lab_UT.scdp.q_RNIABC1D_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u2.q_esr_RNI2EJT_1_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9172\,
            in2 => \_gnd_net_\,
            in3 => \N__9291\,
            lcout => \Lab_UT.scdp.d2eData_1\,
            ltout => \Lab_UT.scdp.d2eData_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.b2a1.lowerTen_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100000"
        )
    port map (
            in0 => \N__9137\,
            in1 => \N__9401\,
            in2 => \N__9160\,
            in3 => \N__9326\,
            lcout => \Lab_UT.scdp.lsBits_6\,
            ltout => \Lab_UT.scdp.lsBits_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lsBitsi.q_esr_1_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9311\,
            in2 => \N__9157\,
            in3 => \N__12356\,
            lcout => \Lab_UT.scdp.lsBitsD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22633\,
            ce => \N__13204\,
            sr => \N__18042\
        );

    \Lab_UT.scdp.lsBitsi.q_esr_3_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__9138\,
            in1 => \N__9402\,
            in2 => \_gnd_net_\,
            in3 => \N__12304\,
            lcout => \Lab_UT.scdp.lsBitsi.lsBitsD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22633\,
            ce => \N__13204\,
            sr => \N__18042\
        );

    \Lab_UT.scdp.lsBitsi.q_esr_6_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100000"
        )
    port map (
            in0 => \N__9403\,
            in1 => \N__9139\,
            in2 => \N__9331\,
            in3 => \N__9315\,
            lcout => \Lab_UT.scdp.lsBitsD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22633\,
            ce => \N__13204\,
            sr => \N__18042\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIO7U41_10_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10824\,
            in1 => \N__10725\,
            in2 => \N__10915\,
            in3 => \N__11779\,
            lcout => \Lab_UT.scdp.d2eData_3_2\,
            ltout => \Lab_UT.scdp.d2eData_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u2.q_esr_RNIEKF71_2_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9346\,
            in3 => \N__9343\,
            lcout => \Lab_UT.scdp.d2eData_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lsBitsi.q_esr_2_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__12357\,
            in1 => \N__9327\,
            in2 => \N__9316\,
            in3 => \N__12305\,
            lcout => \Lab_UT.scdp.lsBitsD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22633\,
            ce => \N__13204\,
            sr => \N__18042\
        );

    \Lab_UT.scdp.pinst0.un12_pValid_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000101000"
        )
    port map (
            in0 => \N__9849\,
            in1 => \N__9292\,
            in2 => \N__14001\,
            in3 => \N__9257\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.pinst0.un12_pValidZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.pinst0.un12_pValid_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9460\,
            in1 => \N__11183\,
            in2 => \N__9277\,
            in3 => \N__9483\,
            lcout => \Lab_UT.scdp.un12_pValid\,
            ltout => \Lab_UT.scdp.un12_pValid_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.pinst0.pValid_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001101110111"
        )
    port map (
            in0 => \N__11184\,
            in1 => \N__9471\,
            in2 => \N__9274\,
            in3 => \N__9234\,
            lcout => \Lab_UT.scdp.pValid_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI9U1R_0_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10768\,
            in1 => \N__10926\,
            in2 => \N__11013\,
            in3 => \N__12544\,
            lcout => \Lab_UT.scdp.d2eData_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNIDHFGA_3_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__9472\,
            in1 => \N__9241\,
            in2 => \_gnd_net_\,
            in3 => \N__9235\,
            lcout => \Lab_UT.scdp.q_RNIDHFGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_esr_RNIDBBI1_2_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9214\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12625\,
            lcout => \Lab_UT.scdp.e2dData_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNITJGS_3_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10949\,
            in1 => \N__11040\,
            in2 => \N__10797\,
            in3 => \N__11160\,
            lcout => \Lab_UT.scdp.N_59_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.pinst0.un12_pValid_1_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000101000"
        )
    port map (
            in0 => \N__9824\,
            in1 => \N__9438\,
            in2 => \N__11848\,
            in3 => \N__9393\,
            lcout => \Lab_UT.scdp.pinst0.un12_pValidZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_RNI239E_4_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12286\,
            in1 => \N__9454\,
            in2 => \_gnd_net_\,
            in3 => \N__18141\,
            lcout => \Lab_UT.scdp.msBitsi.q_esr_RNI239EZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIN7V41_4_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11758\,
            in1 => \N__10980\,
            in2 => \N__10969\,
            in3 => \N__12508\,
            lcout => \Lab_UT.scdp.d2eData_3_4\,
            ltout => \Lab_UT.scdp.d2eData_3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNIIAV0D_0_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11847\,
            in2 => \N__9427\,
            in3 => \N__9374\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.q_RNIIAV0D_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_4_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__17842\,
            in1 => \_gnd_net_\,
            in2 => \N__9424\,
            in3 => \N__9421\,
            lcout => \ufifo.txdataDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNISBU41_3_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10753\,
            in1 => \N__11724\,
            in2 => \N__10900\,
            in3 => \N__10996\,
            lcout => \Lab_UT.scdp.d2eData_3_3\,
            ltout => \Lab_UT.scdp.d2eData_3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_RNIRM8BD_3_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__9375\,
            in1 => \_gnd_net_\,
            in2 => \N__9349\,
            in3 => \N__9825\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.q_RNIRM8BD_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.txdataD_3_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9880\,
            in2 => \N__9871\,
            in3 => \N__17841\,
            lcout => \ufifo.txdataDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_0_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__11869\,
            in1 => \N__14019\,
            in2 => \_gnd_net_\,
            in3 => \N__9848\,
            lcout => \Lab_UT.scdp.byteToDecrypt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22620\,
            ce => 'H',
            sr => \N__18049\
        );

    \Lab_UT.scdp.u1.q_3_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__14020\,
            in1 => \N__11148\,
            in2 => \_gnd_net_\,
            in3 => \N__9826\,
            lcout => \Lab_UT.scdp.byteToDecrypt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22620\,
            ce => 'H',
            sr => \N__18049\
        );

    \ufifo.fifo.wraddr_RNI028U_4_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__9797\,
            in1 => \N__9774\,
            in2 => \N__9744\,
            in3 => \N__9714\,
            lcout => \ufifo.fifo.un1_emptyB_NE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_RNIOP7U_2_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__9680\,
            in1 => \N__9657\,
            in2 => \N__9627\,
            in3 => \N__9597\,
            lcout => OPEN,
            ltout => \ufifo.fifo.un1_emptyB_NE_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.fifo.wraddr_RNIHJBD1_1_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9566\,
            in2 => \N__9547\,
            in3 => \N__9537\,
            lcout => \ufifo.fifo.un1_emptyB_NE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIN78A_0_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__18442\,
            in1 => \N__18953\,
            in2 => \_gnd_net_\,
            in3 => \N__20096\,
            lcout => \Lab_UT.scctrl.g0_16_mb_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_5_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110110000"
        )
    port map (
            in0 => \N__11519\,
            in1 => \N__11301\,
            in2 => \N__11319\,
            in3 => \N__11485\,
            lcout => \ufifo.tx_fsm.cstateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22678\,
            ce => 'H',
            sr => \N__9966\
        );

    \ufifo.tx_fsm.cstate_4_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__9511\,
            in1 => \N__11518\,
            in2 => \_gnd_net_\,
            in3 => \N__12175\,
            lcout => \ufifo.tx_fsm.cstateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22678\,
            ce => 'H',
            sr => \N__9966\
        );

    \buart.Z_tx.bitcount_RNIQOQA1_3_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10134\,
            in1 => \N__10116\,
            in2 => \N__10099\,
            in3 => \N__11964\,
            lcout => \buart__tx_uart_busy_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_1_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100011111000"
        )
    port map (
            in0 => \N__11241\,
            in1 => \N__16069\,
            in2 => \N__10042\,
            in3 => \N__11293\,
            lcout => \ufifo.tx_fsm.cstateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22673\,
            ce => 'H',
            sr => \N__9973\
        );

    \ufifo.fifo.wraddr_RNINV384_1_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10081\,
            in1 => \N__10075\,
            in2 => \N__10066\,
            in3 => \N__10054\,
            lcout => \ufifo.emptyB_0\,
            ltout => \ufifo.emptyB_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNO_0_2_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11517\,
            in2 => \N__10045\,
            in3 => \N__11452\,
            lcout => OPEN,
            ltout => \ufifo.tx_fsm.N_62_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_2_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101000"
        )
    port map (
            in0 => \N__11294\,
            in1 => \N__10038\,
            in2 => \N__10030\,
            in3 => \N__11524\,
            lcout => \ufifo.popFifo\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22673\,
            ce => 'H',
            sr => \N__9973\
        );

    \ufifo.emitcrlf_fsm.cstate_RNO_1_1_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__9943\,
            in1 => \N__11370\,
            in2 => \_gnd_net_\,
            in3 => \N__20283\,
            lcout => \ufifo.emitcrlf_fsm.cstate_srsts_sn_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_7_0_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16163\,
            in1 => \N__17073\,
            in2 => \N__15703\,
            in3 => \N__16960\,
            lcout => \Lab_UT.scctrl.m24_e_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIPVCP_2_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12435\,
            in2 => \_gnd_net_\,
            in3 => \N__10657\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcountlde_i_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__10490\,
            in1 => \N__10552\,
            in2 => \N__9883\,
            in3 => \N__10608\,
            lcout => \buart.Z_rx.N_58\,
            ltout => \buart.Z_rx.N_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_RNIJ3K62_0_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10714\,
            in2 => \N__10222\,
            in3 => \N__10219\,
            lcout => \buart.Z_rx.startbit\,
            ltout => \buart.Z_rx.startbit_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIELQA6_4_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__20787\,
            in1 => \N__10198\,
            in2 => \N__10186\,
            in3 => \N__10183\,
            lcout => \buart.Z_rx.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.g0_17_N_3L3_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__14855\,
            in1 => \N__10486\,
            in2 => \_gnd_net_\,
            in3 => \N__10551\,
            lcout => \Lab_UT.scctrl.g0_17_N_3LZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10603\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10546\,
            in2 => \_gnd_net_\,
            in3 => \N__10147\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12430\,
            in2 => \_gnd_net_\,
            in3 => \N__10144\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10656\,
            in2 => \_gnd_net_\,
            in3 => \N__10141\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_4_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__10357\,
            in1 => \N__10305\,
            in2 => \N__10498\,
            in3 => \N__10138\,
            lcout => \buart__rx_bitcount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22658\,
            ce => \N__10279\,
            sr => \N__18074\
        );

    \buart.Z_rx.bitcount_es_RNIGTPI1_3_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10647\,
            in1 => \N__10589\,
            in2 => \N__10548\,
            in3 => \N__10477\,
            lcout => \buart.Z_rx.bitcount_es_RNIGTPI1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNI4E361_2_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10651\,
            in1 => \N__10534\,
            in2 => \_gnd_net_\,
            in3 => \N__12425\,
            lcout => \buart.Z_rx.N_41_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_3_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__10309\,
            in1 => \N__10360\,
            in2 => \N__10393\,
            in3 => \N__10652\,
            lcout => \buart__rx_bitcount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22653\,
            ce => \N__10278\,
            sr => \N__18069\
        );

    \buart.Z_rx.bitcount_es_1_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000111101100110"
        )
    port map (
            in0 => \N__10547\,
            in1 => \N__10384\,
            in2 => \N__10373\,
            in3 => \N__10307\,
            lcout => \buart__rx_bitcount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22653\,
            ce => \N__10278\,
            sr => \N__18069\
        );

    \buart.Z_rx.bitcount_es_0_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__10306\,
            in1 => \N__10359\,
            in2 => \N__13965\,
            in3 => \N__10590\,
            lcout => \buart__rx_bitcount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22653\,
            ce => \N__10278\,
            sr => \N__18069\
        );

    \buart.Z_rx.bitcount_es_2_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__10358\,
            in1 => \N__10308\,
            in2 => \N__10288\,
            in3 => \N__12426\,
            lcout => \buart__rx_bitcount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22653\,
            ce => \N__10278\,
            sr => \N__18069\
        );

    \Lab_UT.dk.de_bigL_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__10249\,
            in1 => \N__10665\,
            in2 => \N__10258\,
            in3 => \N__10420\,
            lcout => \Lab_UT.de_bigL\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.de_bigL_sx_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__10494\,
            in1 => \N__10535\,
            in2 => \N__14854\,
            in3 => \N__10591\,
            lcout => \Lab_UT.dk.de_bigL_sxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.de_bigL_3_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16549\,
            in1 => \N__16846\,
            in2 => \N__11674\,
            in3 => \N__13474\,
            lcout => \Lab_UT.de_bigL_3\,
            ltout => \Lab_UT.de_bigL_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.g0_17_N_4L5_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__10666\,
            in1 => \N__10243\,
            in2 => \N__10234\,
            in3 => \N__10231\,
            lcout => \Lab_UT.scctrl.g0_17_N_4LZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.de_bigL_0_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17021\,
            in2 => \_gnd_net_\,
            in3 => \N__13250\,
            lcout => \Lab_UT.de_bigL_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_ret_3_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17022\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22646\,
            ce => \N__16753\,
            sr => \N__18075\
        );

    \Lab_UT.dk.de_bigD_1_0_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__16489\,
            in1 => \_gnd_net_\,
            in2 => \N__12434\,
            in3 => \N__10648\,
            lcout => \Lab_UT.dk.de_bigD_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_6_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16854\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22640\,
            ce => \N__16754\,
            sr => \N__18076\
        );

    \Lab_UT.dk.de_bigD_sx_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__10495\,
            in1 => \N__10549\,
            in2 => \N__16899\,
            in3 => \N__10604\,
            lcout => \Lab_UT.dk.de_bigD_sxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIF6D61_4_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__10550\,
            in1 => \N__16853\,
            in2 => \_gnd_net_\,
            in3 => \N__10496\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_es_RNIF6D61Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_fast_RNI639J4_2_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__10444\,
            in1 => \N__10435\,
            in2 => \N__10438\,
            in3 => \N__16433\,
            lcout => \shifter_0_fast_RNI639J4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.de_bigD_0_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16550\,
            in2 => \_gnd_net_\,
            in3 => \N__17019\,
            lcout => \Lab_UT_dk_de_bigD_0\,
            ltout => \Lab_UT_dk_de_bigD_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.de_bigD_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__10429\,
            in1 => \N__16432\,
            in2 => \N__10423\,
            in3 => \N__10419\,
            lcout => \Lab_UT.de_bigD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_7_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10710\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22640\,
            ce => \N__16754\,
            sr => \N__18076\
        );

    \Lab_UT.dk.de_bigE_1_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__17020\,
            in1 => \_gnd_net_\,
            in2 => \N__16900\,
            in3 => \N__16490\,
            lcout => \Lab_UT.dk.de_bigEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_18_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12738\,
            in1 => \N__14893\,
            in2 => \_gnd_net_\,
            in3 => \N__10690\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22634\,
            ce => \N__12469\,
            sr => \N__18078\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_23_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13747\,
            in1 => \N__10839\,
            in2 => \_gnd_net_\,
            in3 => \N__12741\,
            lcout => \Lab_UT.scdp.prng_lfsr_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22634\,
            ce => \N__12469\,
            sr => \N__18078\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_17_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12737\,
            in1 => \N__14929\,
            in2 => \_gnd_net_\,
            in3 => \N__10767\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22634\,
            ce => \N__12469\,
            sr => \N__18078\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_25_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12907\,
            in1 => \N__11014\,
            in2 => \_gnd_net_\,
            in3 => \N__12742\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22634\,
            ce => \N__12469\,
            sr => \N__18078\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_7_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12739\,
            in1 => \N__15412\,
            in2 => \_gnd_net_\,
            in3 => \N__11819\,
            lcout => \Lab_UT.scdp.prng_lfsr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22634\,
            ce => \N__12469\,
            sr => \N__18078\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_14_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13609\,
            in1 => \N__12483\,
            in2 => \_gnd_net_\,
            in3 => \N__12740\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22634\,
            ce => \N__12469\,
            sr => \N__18078\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_15_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12736\,
            in1 => \N__11125\,
            in2 => \_gnd_net_\,
            in3 => \N__10678\,
            lcout => \Lab_UT.scdp.prng_lfsr_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22634\,
            ce => \N__12469\,
            sr => \N__18078\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_30_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13816\,
            in1 => \N__10870\,
            in2 => \_gnd_net_\,
            in3 => \N__12743\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22634\,
            ce => \N__12469\,
            sr => \N__18078\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_22_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12796\,
            in1 => \N__13855\,
            in2 => \_gnd_net_\,
            in3 => \N__10884\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22629\,
            ce => \N__12468\,
            sr => \N__18080\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_19_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13873\,
            in1 => \N__10825\,
            in2 => \_gnd_net_\,
            in3 => \N__12800\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22629\,
            ce => \N__12468\,
            sr => \N__18080\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_10_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12795\,
            in1 => \N__14173\,
            in2 => \_gnd_net_\,
            in3 => \N__10738\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22629\,
            ce => \N__12468\,
            sr => \N__18080\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_4_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15454\,
            in1 => \N__10752\,
            in2 => \_gnd_net_\,
            in3 => \N__12801\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22629\,
            ce => \N__12468\,
            sr => \N__18080\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_26_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__12797\,
            in1 => \_gnd_net_\,
            in2 => \N__13795\,
            in3 => \N__10812\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22629\,
            ce => \N__12468\,
            sr => \N__18080\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_16_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10790\,
            in1 => \N__14947\,
            in2 => \_gnd_net_\,
            in3 => \N__12799\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22629\,
            ce => \N__12468\,
            sr => \N__18080\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_3_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12798\,
            in1 => \N__15052\,
            in2 => \_gnd_net_\,
            in3 => \N__11778\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22629\,
            ce => \N__12468\,
            sr => \N__18080\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_9_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12598\,
            in1 => \N__10927\,
            in2 => \_gnd_net_\,
            in3 => \N__12802\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22629\,
            ce => \N__12468\,
            sr => \N__18080\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_11_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12787\,
            in1 => \N__11107\,
            in2 => \_gnd_net_\,
            in3 => \N__10726\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22626\,
            ce => \N__12466\,
            sr => \N__18082\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_24_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11039\,
            in1 => \N__12450\,
            in2 => \_gnd_net_\,
            in3 => \N__12791\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22626\,
            ce => \N__12466\,
            sr => \N__18082\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_20_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__12788\,
            in1 => \N__10995\,
            in2 => \N__12864\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22626\,
            ce => \N__12466\,
            sr => \N__18082\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_28_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12841\,
            in1 => \N__10899\,
            in2 => \_gnd_net_\,
            in3 => \N__12793\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22626\,
            ce => \N__12466\,
            sr => \N__18082\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_21_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12789\,
            in1 => \N__12577\,
            in2 => \_gnd_net_\,
            in3 => \N__10981\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22626\,
            ce => \N__12466\,
            sr => \N__18082\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_29_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12559\,
            in1 => \N__10968\,
            in2 => \_gnd_net_\,
            in3 => \N__12794\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22626\,
            ce => \N__12466\,
            sr => \N__18082\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_8_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__12790\,
            in1 => \_gnd_net_\,
            in2 => \N__12886\,
            in3 => \N__10950\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22626\,
            ce => \N__12466\,
            sr => \N__18082\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_27_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13699\,
            in1 => \N__10914\,
            in2 => \_gnd_net_\,
            in3 => \N__12792\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22626\,
            ce => \N__12466\,
            sr => \N__18082\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIRBV41_13_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10885\,
            in1 => \N__12484\,
            in2 => \N__10869\,
            in3 => \N__11743\,
            lcout => \Lab_UT.scdp.d2eData_3_5\,
            ltout => \Lab_UT.scdp.d2eData_3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_RNI5V781_1_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11194\,
            in3 => \N__11169\,
            lcout => \Lab_UT.scdp.e2dData_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_1_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__11170\,
            in1 => \N__14040\,
            in2 => \_gnd_net_\,
            in3 => \N__12951\,
            lcout => \Lab_UT.scdp.u0.byteToDecrypt_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22621\,
            ce => 'H',
            sr => \N__18051\
        );

    \Lab_UT.scdp.u0.q_3_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__12952\,
            in1 => \N__11149\,
            in2 => \_gnd_net_\,
            in3 => \N__11161\,
            lcout => \Lab_UT.scdp.u0.byteToDecrypt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22621\,
            ce => 'H',
            sr => \N__18051\
        );

    \Lab_UT.scdp.rxdataD.q_3_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11147\,
            lcout => \Lab_UT.scdp.binValD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22621\,
            ce => 'H',
            sr => \N__18051\
        );

    \Lab_UT.scdp.k1h.q_3_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__11121\,
            in1 => \N__15317\,
            in2 => \N__15249\,
            in3 => \N__13637\,
            lcout => \Lab_UT.scdp.key1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22621\,
            ce => 'H',
            sr => \N__18051\
        );

    \Lab_UT.scdp.k1l.q_3_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__15316\,
            in1 => \N__11106\,
            in2 => \N__15250\,
            in3 => \N__14200\,
            lcout => \Lab_UT.scdp.key1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22621\,
            ce => 'H',
            sr => \N__18051\
        );

    \ufifo.txDataValidD_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__12661\,
            in1 => \N__12634\,
            in2 => \_gnd_net_\,
            in3 => \N__12655\,
            lcout => \ufifo.txDataValidDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22618\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIHLIO_3_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18309\,
            in1 => \N__20155\,
            in2 => \_gnd_net_\,
            in3 => \N__20095\,
            lcout => \Lab_UT.scctrl.g0_14_mb_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNI226B9_4_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100000"
        )
    port map (
            in0 => \N__11225\,
            in1 => \N__11484\,
            in2 => \N__11523\,
            in3 => \N__21011\,
            lcout => OPEN,
            ltout => \ufifo.N_57_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_1_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__11050\,
            in1 => \_gnd_net_\,
            in2 => \N__11044\,
            in3 => \N__11326\,
            lcout => \ufifo.emitcrlf_fsm.cstateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNI7ELR5_4_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11513\,
            in1 => \N__11442\,
            in2 => \_gnd_net_\,
            in3 => \N__16184\,
            lcout => \ufifo.tx_fsm.N_59_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.shifter_ret_3_RNIP72B1_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16297\,
            in1 => \N__16358\,
            in2 => \N__16171\,
            in3 => \N__16956\,
            lcout => \Lab_UT.m61_i_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.g0_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11200\,
            in1 => \N__16162\,
            in2 => \_gnd_net_\,
            in3 => \N__20807\,
            lcout => \Lab_UT.de_bigE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.emitcrlf_fsm.cstate_RNO_0_1_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001100000000"
        )
    port map (
            in0 => \N__11443\,
            in1 => \N__12180\,
            in2 => \N__11385\,
            in3 => \N__20163\,
            lcout => \ufifo.emitcrlf_fsm.cstate_srsts_rn_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNO_0_0_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__11226\,
            in1 => \N__16185\,
            in2 => \_gnd_net_\,
            in3 => \N__21012\,
            lcout => OPEN,
            ltout => \ufifo.tx_fsm.N_72_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_0_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__11320\,
            in1 => \N__11302\,
            in2 => \N__11272\,
            in3 => \N__20164\,
            lcout => \ufifo.cstate_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep2_RNI6VBB5_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22305\,
            in1 => \N__20562\,
            in2 => \N__22093\,
            in3 => \N__17154\,
            lcout => \Lab_UT.scctrl.next_state_1_i_a5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.de_bigE_2_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__16510\,
            in1 => \N__16447\,
            in2 => \N__16971\,
            in3 => \N__17072\,
            lcout => \Lab_UT.dk.de_bigEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_18_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14368\,
            in1 => \N__14433\,
            in2 => \_gnd_net_\,
            in3 => \N__20060\,
            lcout => \Lab_UT.scctrl.g0_i_a7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.state_ret_5_rep2_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22762\,
            lcout => rst_i_3_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIMU571_2_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20563\,
            in1 => \N__23001\,
            in2 => \N__19561\,
            in3 => \N__17502\,
            lcout => \Lab_UT.scctrl.un6_sccDecrypt\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_2_0_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__20786\,
            in1 => \N__11545\,
            in2 => \N__11641\,
            in3 => \N__13017\,
            lcout => \Lab_UT.scctrl.N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.de_cr_0_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16959\,
            in2 => \_gnd_net_\,
            in3 => \N__17066\,
            lcout => OPEN,
            ltout => \Lab_UT.dk.escKey_4_reti_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.shifter_ret_3_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__13433\,
            in1 => \_gnd_net_\,
            in2 => \N__11539\,
            in3 => \N__15665\,
            lcout => \Lab_UT.de_cr_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22650\,
            ce => \N__16757\,
            sr => \N__18077\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_17_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16353\,
            in1 => \N__16958\,
            in2 => \N__16292\,
            in3 => \N__16548\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_i_a3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_14_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010001000100"
        )
    port map (
            in0 => \N__22302\,
            in1 => \N__11536\,
            in2 => \N__11527\,
            in3 => \N__20785\,
            lcout => \Lab_UT.scctrl.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_a9_1_3_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16352\,
            in1 => \N__16155\,
            in2 => \N__16293\,
            in3 => \N__16957\,
            lcout => OPEN,
            ltout => \Lab_UT.g0_i_a9_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_RNIQKK14_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010001000100"
        )
    port map (
            in0 => \N__22303\,
            in1 => \N__16060\,
            in2 => \N__11548\,
            in3 => \N__20784\,
            lcout => \Lab_UT.scctrl.N_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.shifter_ret_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__13374\,
            in1 => \N__11897\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.de_cr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22644\,
            ce => \N__16756\,
            sr => \N__18073\
        );

    \buart.Z_rx.shifter_0_3_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13373\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22644\,
            ce => \N__16756\,
            sr => \N__18073\
        );

    \buart.Z_rx.shifter_0_fast_3_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13375\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart__rx_shifter_0_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22644\,
            ce => \N__16756\,
            sr => \N__18073\
        );

    \buart.Z_rx.shifter_0_0_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15752\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22644\,
            ce => \N__16756\,
            sr => \N__18073\
        );

    \buart.Z_rx.shifter_0_1_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15652\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22644\,
            ce => \N__16756\,
            sr => \N__18073\
        );

    \buart.Z_rx.shifter_0_0_rep1_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15753\,
            lcout => bu_rx_data_0_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22644\,
            ce => \N__16756\,
            sr => \N__18073\
        );

    \buart.Z_rx.shifter_ret_2_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16954\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22644\,
            ce => \N__16756\,
            sr => \N__18073\
        );

    \buart.Z_rx.shifter_0_2_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11898\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22644\,
            ce => \N__16756\,
            sr => \N__18073\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_2_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12419\,
            in2 => \_gnd_net_\,
            in3 => \N__12372\,
            lcout => bu_rx_data_rdy,
            ltout => \bu_rx_data_rdy_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.r1.q_0_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__17810\,
            in1 => \N__11569\,
            in2 => \N__11608\,
            in3 => \N__11563\,
            lcout => \Lab_UT.scctrl.delay1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22638\,
            ce => 'H',
            sr => \N__18041\
        );

    \Lab_UT.scdp.pinst1.un1_pValid_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__13412\,
            in1 => \N__13305\,
            in2 => \_gnd_net_\,
            in3 => \N__16877\,
            lcout => \Lab_UT.un1_pValid\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.r2.q_0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11605\,
            lcout => \Lab_UT.scctrl.delay2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22638\,
            ce => 'H',
            sr => \N__18041\
        );

    \Lab_UT.scctrl.r3.q_0_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11599\,
            lcout => \Lab_UT.scctrl.delay3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22638\,
            ce => 'H',
            sr => \N__18041\
        );

    \Lab_UT.scdp.pinst1.un12_pValid_1_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13357\,
            in1 => \N__16354\,
            in2 => \_gnd_net_\,
            in3 => \N__13411\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.pinst1.un12_pValidZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.pinst1.un7_pValid_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__11586\,
            in1 => \N__16878\,
            in2 => \N__11572\,
            in3 => \N__17059\,
            lcout => \Lab_UT.un7_pValid\,
            ltout => \Lab_UT.un7_pValid_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNIRB726_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__17809\,
            in1 => \N__11562\,
            in2 => \N__11554\,
            in3 => \N__20753\,
            lcout => \Lab_UT.sccEldByte\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_6_RNIFERUH_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__21249\,
            in1 => \N__11713\,
            in2 => \N__21208\,
            in3 => \N__13583\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_1_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_6_RNIL97G01_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010000"
        )
    port map (
            in0 => \N__13584\,
            in1 => \N__18939\,
            in2 => \N__11551\,
            in3 => \N__12786\,
            lcout => \Lab_UT.state_ret_6_RNIL97G01_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_0_sqmuxa_4_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21013\,
            in3 => \N__20209\,
            lcout => \Lab_UT.scctrl.next_state_0_sqmuxa_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.de_bigD_6_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__13252\,
            in1 => \N__11665\,
            in2 => \N__13473\,
            in3 => \N__13509\,
            lcout => \Lab_UT_dk_de_bigD_6\,
            ltout => \Lab_UT_dk_de_bigD_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.de_bigE_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16136\,
            in1 => \N__11707\,
            in2 => \N__11701\,
            in3 => \N__20719\,
            lcout => \Lab_UT.de_bigE\,
            ltout => \Lab_UT.de_bigE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_6_RNIJMNGE_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__13528\,
            in1 => \N__17135\,
            in2 => \N__11698\,
            in3 => \N__17198\,
            lcout => \Lab_UT.scctrl.next_state_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.val_i_0_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101111110010"
        )
    port map (
            in0 => \N__14867\,
            in1 => \N__15680\,
            in2 => \N__11689\,
            in3 => \N__16146\,
            lcout => \Lab_UT.scdp.N_39\,
            ltout => \Lab_UT.scdp.N_39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.rxdataD.q_0_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11695\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.scdp.binValD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22628\,
            ce => 'H',
            sr => \N__18046\
        );

    \Lab_UT.scdp.a2b.val_0_o2_3_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__16879\,
            in1 => \N__13469\,
            in2 => \N__13324\,
            in3 => \N__11679\,
            lcout => \Lab_UT.scdp.a2b.N_50\,
            ltout => \Lab_UT.scdp.a2b.N_50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.val_i_o2_0_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11692\,
            in3 => \N__11932\,
            lcout => \Lab_UT.scdp.a2b.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_8_0_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14866\,
            in1 => \N__13468\,
            in2 => \N__11935\,
            in3 => \N__11678\,
            lcout => \Lab_UT.scctrl.m24_e_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.val_i_o2_1_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__11619\,
            in1 => \N__11933\,
            in2 => \_gnd_net_\,
            in3 => \N__16142\,
            lcout => \Lab_UT.scdp.a2b.N_53\,
            ltout => \Lab_UT.scdp.a2b.N_53_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.val_i_1_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__14868\,
            in1 => \N__15758\,
            in2 => \N__11872\,
            in3 => \N__15681\,
            lcout => \Lab_UT.scdp.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_0_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__11865\,
            in1 => \N__11838\,
            in2 => \_gnd_net_\,
            in3 => \N__12945\,
            lcout => \Lab_UT.scdp.byteToDecrypt_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22628\,
            ce => 'H',
            sr => \N__18046\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_6_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11742\,
            in1 => \N__15529\,
            in2 => \_gnd_net_\,
            in3 => \N__12751\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22624\,
            ce => \N__12467\,
            sr => \N__18083\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_RNO_0_0_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12500\,
            in1 => \N__11741\,
            in2 => \N__11823\,
            in3 => \N__11777\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.lfsrInst.prng_lfsr_next_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__13680\,
            in1 => \N__11796\,
            in2 => \N__11782\,
            in3 => \N__12748\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22624\,
            ce => \N__12467\,
            sr => \N__18083\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_2_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12747\,
            in1 => \N__13665\,
            in2 => \_gnd_net_\,
            in3 => \N__12522\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22624\,
            ce => \N__12467\,
            sr => \N__18083\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_5_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15838\,
            in1 => \N__11757\,
            in2 => \_gnd_net_\,
            in3 => \N__12750\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22624\,
            ce => \N__12467\,
            sr => \N__18083\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_12_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12745\,
            in1 => \N__13654\,
            in2 => \_gnd_net_\,
            in3 => \N__11725\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22624\,
            ce => \N__12467\,
            sr => \N__18083\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_1_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15343\,
            in1 => \N__12540\,
            in2 => \_gnd_net_\,
            in3 => \N__12749\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22624\,
            ce => \N__12467\,
            sr => \N__18083\
        );

    \Lab_UT.scdp.lfsrInst.prng_lfsr_13_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__12746\,
            in1 => \_gnd_net_\,
            in2 => \N__12507\,
            in3 => \N__12613\,
            lcout => \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22624\,
            ce => \N__12467\,
            sr => \N__18083\
        );

    \Lab_UT.scdp.k3l.q_0_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__15497\,
            in1 => \N__12451\,
            in2 => \N__15272\,
            in3 => \N__13722\,
            lcout => \Lab_UT.scdp.key3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => 'H',
            sr => \N__18052\
        );

    \Lab_UT.scdp.rddataDV.q_0_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12439\,
            in2 => \_gnd_net_\,
            in3 => \N__12379\,
            lcout => \Lab_UT.scdp.binVal_ValidD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => 'H',
            sr => \N__18052\
        );

    \Lab_UT.scdp.lsBitsi.q_0_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__13181\,
            in1 => \N__12361\,
            in2 => \N__12333\,
            in3 => \N__12313\,
            lcout => \Lab_UT.scdp.lsBitsD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => 'H',
            sr => \N__18052\
        );

    \Lab_UT.scdp.lsBitsi.q_4_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__12285\,
            in1 => \N__12312\,
            in2 => \_gnd_net_\,
            in3 => \N__13183\,
            lcout => \Lab_UT.scdp.lsBitsD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => 'H',
            sr => \N__18052\
        );

    \Lab_UT.scdp.msBitsi.q_3_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__13182\,
            in1 => \N__12268\,
            in2 => \N__12207\,
            in3 => \N__12229\,
            lcout => \Lab_UT.scdp.msBitsD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => 'H',
            sr => \N__18052\
        );

    \buart.Z_tx.bitcount_0_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110101000000000"
        )
    port map (
            in0 => \N__11960\,
            in1 => \N__12184\,
            in2 => \N__12115\,
            in3 => \N__12052\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => 'H',
            sr => \N__18052\
        );

    \Lab_UT.scctrl.state_ret_13_RNIQ72741_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13638\,
            in1 => \N__15034\,
            in2 => \_gnd_net_\,
            in3 => \N__14983\,
            lcout => \Lab_UT.state_ret_13_RNIQ72741_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.r4.q_0_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12654\,
            lcout => \Lab_UT.scctrl.r4.delay4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => 'H',
            sr => \N__18052\
        );

    \Lab_UT.scdp.u1.q_esr_2_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__15682\,
            in1 => \N__15776\,
            in2 => \_gnd_net_\,
            in3 => \N__15809\,
            lcout => \Lab_UT.scdp.u1.byteToDecrypt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22617\,
            ce => \N__14047\,
            sr => \N__18054\
        );

    \Lab_UT.scctrl.state_2_RNI44QH41_2_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13771\,
            in1 => \N__18199\,
            in2 => \_gnd_net_\,
            in3 => \N__14984\,
            lcout => \Lab_UT.state_2_RNI44QH41_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNI416G41_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14986\,
            in1 => \N__14676\,
            in2 => \_gnd_net_\,
            in3 => \N__13837\,
            lcout => \Lab_UT.state_ret_14_RNI416G41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIF0RJ41_2_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13726\,
            in1 => \N__18220\,
            in2 => \_gnd_net_\,
            in3 => \N__14985\,
            lcout => \Lab_UT.state_2_RNIF0RJ41_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.k1h.q_1_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__12612\,
            in1 => \N__15384\,
            in2 => \N__15274\,
            in3 => \N__13639\,
            lcout => \Lab_UT.scdp.key1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22615\,
            ce => 'H',
            sr => \N__18055\
        );

    \Lab_UT.scdp.k1l.q_1_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__15383\,
            in1 => \N__15231\,
            in2 => \N__12597\,
            in3 => \N__14199\,
            lcout => \Lab_UT.scdp.key1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22615\,
            ce => 'H',
            sr => \N__18055\
        );

    \Lab_UT.scdp.k2h.q_1_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__12573\,
            in1 => \N__15385\,
            in2 => \N__15275\,
            in3 => \N__13768\,
            lcout => \Lab_UT.scdp.key2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22615\,
            ce => 'H',
            sr => \N__18055\
        );

    \Lab_UT.scdp.k3h.q_1_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__13835\,
            in1 => \N__15233\,
            in2 => \N__15391\,
            in3 => \N__12558\,
            lcout => \Lab_UT.scdp.key3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22615\,
            ce => 'H',
            sr => \N__18055\
        );

    \Lab_UT.scdp.k3l.q_1_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__15229\,
            in1 => \N__15386\,
            in2 => \N__12906\,
            in3 => \N__13723\,
            lcout => \Lab_UT.scdp.key3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22615\,
            ce => 'H',
            sr => \N__18055\
        );

    \Lab_UT.scdp.k1l.q_0_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__15498\,
            in1 => \N__15230\,
            in2 => \N__12885\,
            in3 => \N__14198\,
            lcout => \Lab_UT.scdp.key1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22615\,
            ce => 'H',
            sr => \N__18055\
        );

    \Lab_UT.scdp.k2h.q_0_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__15228\,
            in1 => \N__15499\,
            in2 => \N__12865\,
            in3 => \N__13767\,
            lcout => \Lab_UT.scdp.key2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22615\,
            ce => 'H',
            sr => \N__18055\
        );

    \Lab_UT.scdp.k3h.q_0_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__13834\,
            in1 => \N__15232\,
            in2 => \N__15509\,
            in3 => \N__12837\,
            lcout => \Lab_UT.scdp.key3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22615\,
            ce => 'H',
            sr => \N__18055\
        );

    \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_i_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__12819\,
            in1 => \N__14117\,
            in2 => \N__14155\,
            in3 => \N__12744\,
            lcout => \Lab_UT.scdp.lfsrInst.un1_ldLFSR_1_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNIMEE3_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22268\,
            in1 => \N__19698\,
            in2 => \_gnd_net_\,
            in3 => \N__21955\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.un1_state_inv_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_12_RNIUQFK_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101110000"
        )
    port map (
            in0 => \N__20256\,
            in1 => \N__20577\,
            in2 => \N__12670\,
            in3 => \N__18955\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.state_ret_12_RNIUQFKZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_12_RNIMJCP8_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001110"
        )
    port map (
            in0 => \N__13048\,
            in1 => \N__14118\,
            in2 => \N__12667\,
            in3 => \N__19150\,
            lcout => \Lab_UT.state_ret_12_RNIMJCP8_0\,
            ltout => \Lab_UT.state_ret_12_RNIMJCP8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.r5.q_0_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12664\,
            in3 => \N__14153\,
            lcout => \Lab_UT.scctrl.delayload\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22614\,
            ce => 'H',
            sr => \N__18058\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_5_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__19699\,
            in1 => \N__20576\,
            in2 => \_gnd_net_\,
            in3 => \N__22269\,
            lcout => \Lab_UT.scctrl.g0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNIM6P13_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__21127\,
            in1 => \N__17623\,
            in2 => \_gnd_net_\,
            in3 => \N__21014\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNISBDB3_2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__20084\,
            in1 => \_gnd_net_\,
            in2 => \N__12922\,
            in3 => \N__20308\,
            lcout => \Lab_UT.scctrl.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNINMBN3_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__20083\,
            in1 => \N__19695\,
            in2 => \N__13495\,
            in3 => \N__20803\,
            lcout => \Lab_UT.scctrl.g0_i_a9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNI07T4_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19696\,
            in1 => \N__20082\,
            in2 => \N__22339\,
            in3 => \N__20462\,
            lcout => \Lab_UT.scctrl.G_23_0_a9_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNI4DGV4_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__14206\,
            in1 => \N__13552\,
            in2 => \N__16408\,
            in3 => \N__20804\,
            lcout => \Lab_UT.scctrl.g0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.state_ret_5_rep1_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22768\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rst_i_3_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22679\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIO386G1_2_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__14473\,
            in1 => \N__14346\,
            in2 => \_gnd_net_\,
            in3 => \N__14331\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.un1_state_3_1_reti_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_10_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010101010101"
        )
    port map (
            in0 => \N__22767\,
            in1 => \N__14212\,
            in2 => \N__12919\,
            in3 => \N__14290\,
            lcout => \Lab_UT.scctrl.state_retZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22679\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNI0D9CA_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__18947\,
            in1 => \N__20076\,
            in2 => \N__12916\,
            in3 => \N__13021\,
            lcout => \Lab_UT.scctrl.g0_16_mb_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.state_ret_5_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22780\,
            lcout => rst_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_11_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21424\,
            in1 => \N__20075\,
            in2 => \N__21782\,
            in3 => \N__22090\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_4_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__12994\,
            in1 => \N__19425\,
            in2 => \N__12985\,
            in3 => \N__21006\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12961\,
            in1 => \N__12976\,
            in2 => \N__12982\,
            in3 => \N__18967\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_0_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__12970\,
            in1 => \N__14289\,
            in2 => \N__12979\,
            in3 => \N__14521\,
            lcout => \Lab_UT.scctrl.N_1_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_6_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__20077\,
            in1 => \N__23021\,
            in2 => \N__21439\,
            in3 => \N__19166\,
            lcout => \Lab_UT.scctrl.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_2_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20331\,
            in2 => \N__20097\,
            in3 => \N__17888\,
            lcout => \Lab_UT.scctrl.g2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_7_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__21007\,
            in1 => \_gnd_net_\,
            in2 => \N__21173\,
            in3 => \N__20071\,
            lcout => \Lab_UT.scctrl.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_10_RNIPCFBB_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000001"
        )
    port map (
            in0 => \N__13110\,
            in1 => \N__14146\,
            in2 => \N__13096\,
            in3 => \N__13059\,
            lcout => \Lab_UT.sccDnibble1En\,
            ltout => \Lab_UT.sccDnibble1En_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u0.q_esr_RNO_2_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13129\,
            in3 => \N__14087\,
            lcout => \Lab_UT.scdp.u0.sccDnibble1En_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_RNI658G_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21742\,
            in1 => \N__17554\,
            in2 => \N__21440\,
            in3 => \N__21927\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_1_sqmuxa_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_RNI4CFD9_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__18612\,
            in1 => \_gnd_net_\,
            in2 => \N__13114\,
            in3 => \N__18771\,
            lcout => \Lab_UT.scctrl.next_state_1_sqmuxa_3\,
            ltout => \Lab_UT.scctrl.next_state_1_sqmuxa_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__13111\,
            in1 => \N__22781\,
            in2 => \N__13099\,
            in3 => \N__13095\,
            lcout => \Lab_UT.scctrl.nibbleInZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22666\,
            ce => \N__13081\,
            sr => \N__13066\
        );

    \Lab_UT.scctrl.state_ret_8_RNIQ79K1_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__13044\,
            in1 => \N__21950\,
            in2 => \N__21791\,
            in3 => \N__21428\,
            lcout => \Lab_UT.sccDecrypt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_11_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__21743\,
            in1 => \N__18611\,
            in2 => \N__14278\,
            in3 => \N__18763\,
            lcout => \Lab_UT.scctrl.N_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_RNIJLL09_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__18764\,
            in1 => \N__15985\,
            in2 => \N__18627\,
            in3 => \N__21949\,
            lcout => \Lab_UT.scctrl.N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNIHB2UD_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000111111"
        )
    port map (
            in0 => \N__13030\,
            in1 => \N__20928\,
            in2 => \N__14269\,
            in3 => \N__13016\,
            lcout => \Lab_UT.next_state_rst_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNIK9603_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010000"
        )
    port map (
            in0 => \N__18913\,
            in1 => \N__20927\,
            in2 => \N__17840\,
            in3 => \N__13000\,
            lcout => \Lab_UT.scctrl.EmsLoaded\,
            ltout => \Lab_UT.scctrl.EmsLoaded_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNIEOE1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13210\,
            in3 => \N__17829\,
            lcout => \Lab_UT.sccElsBitsLd\,
            ltout => \Lab_UT.sccElsBitsLd_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.msBitsi.q_esr_ctle_6_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13207\,
            in3 => \N__14094\,
            lcout => \Lab_UT.scdp.sccElsBitsLd_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNO_6_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18914\,
            in1 => \N__20184\,
            in2 => \_gnd_net_\,
            in3 => \N__20078\,
            lcout => \Lab_UT.scctrl.G_24_i_a4_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.lsBitsi.q_5_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13146\,
            in2 => \_gnd_net_\,
            in3 => \N__13170\,
            lcout => \Lab_UT.scdp.lsBitsi.lsBitsD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22659\,
            ce => 'H',
            sr => \N__18044\
        );

    \Lab_UT.dk.shifter_ret_3_RNIA82U_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__16270\,
            in1 => \N__16341\,
            in2 => \_gnd_net_\,
            in3 => \N__16944\,
            lcout => \Lab_UT_dk_de_cr_12_1\,
            ltout => \Lab_UT_dk_de_cr_12_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.shifter_ret_3_RNIJC3U2_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16546\,
            in2 => \N__13135\,
            in3 => \N__20718\,
            lcout => \L4_PrintBuf\,
            ltout => \L4_PrintBuf_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep1_RNIHA8U3_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110101"
        )
    port map (
            in0 => \N__17576\,
            in1 => \_gnd_net_\,
            in2 => \N__13132\,
            in3 => \N__14701\,
            lcout => \Lab_UT.state_ret_8_rep1_RNIHA8U3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI5GLD_0_3_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20521\,
            in2 => \_gnd_net_\,
            in3 => \N__17499\,
            lcout => \Lab_UT.scctrl.g0_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.g1_i_a7_2_3_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16547\,
            in1 => \N__16342\,
            in2 => \N__16291\,
            in3 => \N__16945\,
            lcout => \Lab_UT.scctrl.g1_i_a7_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_8_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__20911\,
            in1 => \N__20018\,
            in2 => \N__21200\,
            in3 => \N__13264\,
            lcout => \Lab_UT.scctrl.g0_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI6J7KA_3_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__17500\,
            in1 => \N__19069\,
            in2 => \N__23073\,
            in3 => \N__20910\,
            lcout => \Lab_UT.N_190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g1_1_o2_0_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__20912\,
            in1 => \N__14404\,
            in2 => \N__19118\,
            in3 => \N__13519\,
            lcout => \Lab_UT.scdp.a2b.g1_1_o2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_fast_0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15754\,
            lcout => bu_rx_data_fast_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22647\,
            ce => \N__16755\,
            sr => \N__18079\
        );

    \Lab_UT.dk.un7_de_hex_x0_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000010011"
        )
    port map (
            in0 => \N__16500\,
            in1 => \N__13216\,
            in2 => \N__13510\,
            in3 => \N__13258\,
            lcout => OPEN,
            ltout => \Lab_UT.dk.un7_de_hex_xZ0Z0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.un7_de_hex_ns_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__13251\,
            in1 => \_gnd_net_\,
            in2 => \N__13231\,
            in3 => \N__13964\,
            lcout => \Lab_UT.dk.un7_de_hex_0\,
            ltout => \Lab_UT.dk.un7_de_hex_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.de_hex_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101110111"
        )
    port map (
            in0 => \N__13278\,
            in1 => \N__20713\,
            in2 => \N__13228\,
            in3 => \N__13483\,
            lcout => \Lab_UT.de_hex_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.un4_de_hex_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100000"
        )
    port map (
            in0 => \N__13482\,
            in1 => \N__13225\,
            in2 => \N__20757\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.un4_de_hex\,
            ltout => \Lab_UT.un4_de_hex_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNI68R1A_2_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__20752\,
            in1 => \N__14359\,
            in2 => \N__13219\,
            in3 => \N__13279\,
            lcout => \Lab_UT.N_191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_fast_1_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15651\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart__rx_shifter_0_fast_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22647\,
            ce => \N__16755\,
            sr => \N__18079\
        );

    \buart.Z_rx.shifter_ret_1_fast_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15650\,
            lcout => \buart__rx_shifter_ret_1_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22647\,
            ce => \N__16755\,
            sr => \N__18079\
        );

    \Lab_UT.scctrl.g0_i_o9_0_2_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__13408\,
            in1 => \N__13350\,
            in2 => \N__13323\,
            in3 => \N__16890\,
            lcout => \Lab_UT.scctrl.g0_i_o9_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_4_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13410\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22641\,
            ce => \N__16758\,
            sr => \N__18081\
        );

    \buart.Z_rx.shifter_0_5_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17049\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22641\,
            ce => \N__16758\,
            sr => \N__18081\
        );

    \Lab_UT.dk.un4_de_hex_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17048\,
            in1 => \N__13406\,
            in2 => \N__16940\,
            in3 => \N__13464\,
            lcout => \Lab_UT.dk.un4_de_hexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_ret_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__13409\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22641\,
            ce => \N__16758\,
            sr => \N__18081\
        );

    \Lab_UT.dk.un1_de_hex_2_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13407\,
            in1 => \N__13349\,
            in2 => \N__13322\,
            in3 => \N__16886\,
            lcout => \Lab_UT.un1_de_hex_2\,
            ltout => \Lab_UT.un1_de_hex_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.un1_de_hex_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13267\,
            in3 => \N__20717\,
            lcout => \Lab_UT.un1_de_hex\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_fast_RNI55RL_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__16941\,
            in1 => \N__19915\,
            in2 => \N__14443\,
            in3 => \N__19211\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_i_a9_3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_fast_RNI86TJ1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16164\,
            in1 => \N__16305\,
            in2 => \N__13555\,
            in3 => \N__16367\,
            lcout => \Lab_UT.scctrl.g0_i_a9_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNO_9_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__16942\,
            in1 => \N__16165\,
            in2 => \N__16372\,
            in3 => \N__16306\,
            lcout => \Lab_UT.scctrl.m26_i_o4_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_fast_RNI7JDJ_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19212\,
            in1 => \N__14442\,
            in2 => \_gnd_net_\,
            in3 => \N__21673\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_1_0_a5_2_out_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_fast_RNI21I2A_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010101"
        )
    port map (
            in0 => \N__13915\,
            in1 => \N__18591\,
            in2 => \N__13537\,
            in3 => \N__18730\,
            lcout => \Lab_UT.next_state_1_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_0_1_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19916\,
            in1 => \N__17686\,
            in2 => \_gnd_net_\,
            in3 => \N__14622\,
            lcout => \Lab_UT.state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22635\,
            ce => 'H',
            sr => \N__18048\
        );

    \Lab_UT.scctrl.state_ret_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__14623\,
            in1 => \N__17687\,
            in2 => \N__14482\,
            in3 => \N__19917\,
            lcout => \Lab_UT.scctrl.N_222_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22635\,
            ce => 'H',
            sr => \N__18048\
        );

    \Lab_UT.scctrl.state_ret_RNILUJH_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19662\,
            in1 => \N__21941\,
            in2 => \_gnd_net_\,
            in3 => \N__13534\,
            lcout => \Lab_UT.scctrl.next_state76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_6_RNICI45_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21426\,
            in1 => \N__21248\,
            in2 => \_gnd_net_\,
            in3 => \N__17343\,
            lcout => \Lab_UT.scctrl.next_state_3_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g1_1_a3_0_0_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__21427\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23088\,
            lcout => \Lab_UT.scdp.a2b.g1_1_a3_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.k0l.q_0_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__15489\,
            in1 => \N__13681\,
            in2 => \N__15276\,
            in3 => \N__15075\,
            lcout => \Lab_UT.scdp.key0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22630\,
            ce => 'H',
            sr => \N__18053\
        );

    \Lab_UT.scdp.k0l.q_2_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__15076\,
            in1 => \N__15240\,
            in2 => \N__13669\,
            in3 => \N__15567\,
            lcout => \Lab_UT.scdp.key0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22630\,
            ce => 'H',
            sr => \N__18053\
        );

    \Lab_UT.scdp.k1h.q_0_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__15490\,
            in1 => \N__13653\,
            in2 => \N__15277\,
            in3 => \N__13636\,
            lcout => \Lab_UT.scdp.key1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22630\,
            ce => 'H',
            sr => \N__18053\
        );

    \Lab_UT.scdp.k1h.q_2_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__13635\,
            in1 => \N__13602\,
            in2 => \N__15286\,
            in3 => \N__15568\,
            lcout => \Lab_UT.scdp.key1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22630\,
            ce => 'H',
            sr => \N__18053\
        );

    \Lab_UT.scctrl.state_0_RNIBE791_1_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21698\,
            in2 => \N__23094\,
            in3 => \N__13911\,
            lcout => \Lab_UT.scctrl.next_state77\,
            ltout => \Lab_UT.scctrl.next_state77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_3_RNIHF1E3_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13884\,
            in1 => \N__14727\,
            in2 => \N__13588\,
            in3 => \N__14995\,
            lcout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNIG62DM_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__15030\,
            in1 => \N__19108\,
            in2 => \N__20222\,
            in3 => \N__13585\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNI91DN31_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101001111"
        )
    port map (
            in0 => \N__19109\,
            in1 => \N__20188\,
            in2 => \N__13567\,
            in3 => \N__13894\,
            lcout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i\,
            ltout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_0_RNIKFK051_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13564\,
            in2 => \N__13558\,
            in3 => \N__15081\,
            lcout => \Lab_UT.state_0_RNIKFK051_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep1_RNIT6TH_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19210\,
            in2 => \_gnd_net_\,
            in3 => \N__17440\,
            lcout => \Lab_UT.scctrl.next_state77_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIDHLT5_2_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__18198\,
            in1 => \N__18216\,
            in2 => \N__14677\,
            in3 => \N__13900\,
            lcout => \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_1_0_tz_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_RNIUV0941_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__15433\,
            in1 => \_gnd_net_\,
            in2 => \N__13888\,
            in3 => \N__14982\,
            lcout => \Lab_UT.state_ret_RNIUV0941_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.k2l.q_3_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__13869\,
            in1 => \N__15322\,
            in2 => \N__15251\,
            in3 => \N__14911\,
            lcout => \Lab_UT.scdp.key2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22622\,
            ce => 'H',
            sr => \N__18056\
        );

    \Lab_UT.scdp.k2h.q_2_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__13851\,
            in1 => \N__15558\,
            in2 => \N__15247\,
            in3 => \N__13769\,
            lcout => \Lab_UT.scdp.key2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22622\,
            ce => 'H',
            sr => \N__18056\
        );

    \Lab_UT.scdp.k3h.q_2_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__15559\,
            in1 => \N__15184\,
            in2 => \N__13815\,
            in3 => \N__13836\,
            lcout => \Lab_UT.scdp.key3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22622\,
            ce => 'H',
            sr => \N__18056\
        );

    \Lab_UT.scdp.k3l.q_2_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__15183\,
            in1 => \N__15560\,
            in2 => \N__13791\,
            in3 => \N__13724\,
            lcout => \Lab_UT.scdp.key3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22622\,
            ce => 'H',
            sr => \N__18056\
        );

    \Lab_UT.scdp.k2h.q_3_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__13770\,
            in1 => \N__13740\,
            in2 => \N__15252\,
            in3 => \N__15323\,
            lcout => \Lab_UT.scdp.key2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22622\,
            ce => 'H',
            sr => \N__18056\
        );

    \Lab_UT.scdp.k3l.q_3_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__15321\,
            in1 => \N__13695\,
            in2 => \N__15248\,
            in3 => \N__13725\,
            lcout => \Lab_UT.scdp.key3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22622\,
            ce => 'H',
            sr => \N__18056\
        );

    \Lab_UT.scctrl.state_ret_13_RNIHUNI41_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14194\,
            in1 => \N__14731\,
            in2 => \_gnd_net_\,
            in3 => \N__14980\,
            lcout => \Lab_UT.state_ret_13_RNIHUNI41_0\,
            ltout => \Lab_UT.state_ret_13_RNIHUNI41_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.k1l.q_2_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__15182\,
            in1 => \N__15557\,
            in2 => \N__14176\,
            in3 => \N__14169\,
            lcout => \Lab_UT.scdp.key1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22622\,
            ce => 'H',
            sr => \N__18056\
        );

    \Lab_UT.scctrl.state_ret_8_RNIQ79K1_0_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14154\,
            in2 => \_gnd_net_\,
            in3 => \N__14119\,
            lcout => \Lab_UT.sccDnibble2En\,
            ltout => \Lab_UT.sccDnibble2En_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_esr_RNO_2_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14104\,
            in3 => \N__14101\,
            lcout => \Lab_UT.scdp.u1.sccDnibble2En_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.u1.q_1_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__14041\,
            in1 => \N__13988\,
            in2 => \_gnd_net_\,
            in3 => \N__14013\,
            lcout => \Lab_UT.scdp.byteToDecrypt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22616\,
            ce => 'H',
            sr => \N__18060\
        );

    \Lab_UT.scctrl.next_state_2_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13963\,
            lcout => \Lab_UT.scctrl.next_state_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22695\,
            ce => \N__14792\,
            sr => \N__18087\
        );

    \Lab_UT.scctrl.state_2_RNICEINI_2_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__14218\,
            in1 => \N__18621\,
            in2 => \N__14233\,
            in3 => \N__18781\,
            lcout => \Lab_UT.scctrl.G_23_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIGC1Q_2_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20081\,
            in1 => \N__19555\,
            in2 => \_gnd_net_\,
            in3 => \N__23065\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_i_a9_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_RNI7NLQ7_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__19163\,
            in1 => \N__20463\,
            in2 => \N__13918\,
            in3 => \N__22335\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_RNIK1DPL_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__18623\,
            in1 => \N__14248\,
            in2 => \N__14242\,
            in3 => \N__14239\,
            lcout => \Lab_UT.scctrl.g0_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIU7GR_2_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__19556\,
            in1 => \N__17497\,
            in2 => \N__20512\,
            in3 => \N__20079\,
            lcout => \Lab_UT.scctrl.G_23_0_a9_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_10_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__20080\,
            in1 => \N__22334\,
            in2 => \N__22065\,
            in3 => \N__20458\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_i_a10_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_8_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18622\,
            in2 => \N__14221\,
            in3 => \N__18782\,
            lcout => \Lab_UT.scctrl.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNIGVQU8_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__16003\,
            in1 => \N__20593\,
            in2 => \N__15997\,
            in3 => \N__19162\,
            lcout => \Lab_UT.scctrl.G_23_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNIK9N021_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__15914\,
            in1 => \N__15856\,
            in2 => \N__15897\,
            in3 => \N__15943\,
            lcout => \Lab_UT.scctrl.N_2ctr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNIRRFK_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110110011"
        )
    port map (
            in0 => \N__20091\,
            in1 => \N__17336\,
            in2 => \N__22422\,
            in3 => \N__21764\,
            lcout => \Lab_UT.scctrl.g0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_12_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__14302\,
            in1 => \N__14311\,
            in2 => \N__17095\,
            in3 => \N__14317\,
            lcout => \Lab_UT.state_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_9_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101011111"
        )
    port map (
            in0 => \N__20089\,
            in1 => \N__21419\,
            in2 => \N__21172\,
            in3 => \N__21762\,
            lcout => \Lab_UT.scctrl.g0_i_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__14475\,
            in1 => \N__14347\,
            in2 => \_gnd_net_\,
            in3 => \N__14335\,
            lcout => \Lab_UT.un1_state_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep2_RNIR10T_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20090\,
            in1 => \N__21420\,
            in2 => \N__22091\,
            in3 => \N__21763\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_23_0_a9_4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNIEA5S3_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__21126\,
            in1 => \N__20092\,
            in2 => \N__14320\,
            in3 => \N__21023\,
            lcout => \Lab_UT.scctrl.G_23_0_3\,
            ltout => \Lab_UT.scctrl.G_23_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNIDDIN51_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__14310\,
            in1 => \N__14301\,
            in2 => \N__14293\,
            in3 => \N__17091\,
            lcout => \Lab_UT.scctrl.N_3ctr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_16_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20088\,
            in2 => \_gnd_net_\,
            in3 => \N__19237\,
            lcout => \Lab_UT.scctrl.g0_i_a7_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_RNILGT2_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22312\,
            in2 => \_gnd_net_\,
            in3 => \N__20443\,
            lcout => \Lab_UT.scctrl.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNIGKQK_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20442\,
            in1 => \N__22414\,
            in2 => \N__22333\,
            in3 => \N__23020\,
            lcout => \Lab_UT.scctrl.next_state_1_i_a5_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep1_RNIS10T_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__19293\,
            in1 => \N__21376\,
            in2 => \N__21128\,
            in3 => \N__21760\,
            lcout => \Lab_UT.scctrl.N_166_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_RNI7UQVB_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__21869\,
            in1 => \N__14254\,
            in2 => \N__21202\,
            in3 => \N__20988\,
            lcout => \Lab_UT.scctrl.g0_0_i_2\,
            ltout => \Lab_UT.scctrl.g0_0_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_fast_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__15896\,
            in1 => \N__15922\,
            in2 => \N__14446\,
            in3 => \N__15859\,
            lcout => \Lab_UT.scctrl.state_i_3_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_6_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000100000"
        )
    port map (
            in0 => \N__21868\,
            in1 => \N__14410\,
            in2 => \N__21201\,
            in3 => \N__20987\,
            lcout => \Lab_UT.scctrl.g0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g1_1_o3_1_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__21377\,
            in1 => \N__21867\,
            in2 => \N__21129\,
            in3 => \N__21761\,
            lcout => \Lab_UT.scdp.a2b.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_0_RNI2GENA_1_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__21768\,
            in1 => \N__18599\,
            in2 => \N__16417\,
            in3 => \N__18772\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNI8MD1N_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__14392\,
            in1 => \N__16009\,
            in2 => \N__14377\,
            in3 => \N__14374\,
            lcout => \Lab_UT.next_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep1_RNIP54M_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20062\,
            in1 => \N__19310\,
            in2 => \_gnd_net_\,
            in3 => \N__19238\,
            lcout => \Lab_UT.scctrl.G_21_i_a7_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep2_RNIT10T_0_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__21767\,
            in1 => \N__21161\,
            in2 => \N__22101\,
            in3 => \N__21401\,
            lcout => \Lab_UT.N_166_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI6J7KA_0_3_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__17482\,
            in1 => \N__19147\,
            in2 => \N__23064\,
            in3 => \N__20989\,
            lcout => \Lab_UT.scctrl.N_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_fast_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20630\,
            lcout => \Lab_UT.scctrl.state_i_3_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNI81K41_2_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19537\,
            in1 => \N__21765\,
            in2 => \_gnd_net_\,
            in3 => \N__22993\,
            lcout => \Lab_UT.scctrl.next_state_1_0_a5_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep2_RNIT10T_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__21766\,
            in1 => \N__21160\,
            in2 => \N__22100\,
            in3 => \N__21400\,
            lcout => \Lab_UT.scctrl.N_166_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.state_ret_5_rep2_RNIKU94_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__17616\,
            in1 => \N__18918\,
            in2 => \_gnd_net_\,
            in3 => \N__20051\,
            lcout => OPEN,
            ltout => \N_127_i_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNI2UI47_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__20930\,
            in1 => \N__21165\,
            in2 => \N__14509\,
            in3 => \N__14506\,
            lcout => \Lab_UT.scctrl.N_127_i_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_4_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__18355\,
            in1 => \N__16237\,
            in2 => \N__21195\,
            in3 => \N__20929\,
            lcout => \Lab_UT.scdp.a2b.g0_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g1_i_a4_0_2_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000000000"
        )
    port map (
            in0 => \N__20931\,
            in1 => \N__14497\,
            in2 => \N__17626\,
            in3 => \N__16669\,
            lcout => OPEN,
            ltout => \Lab_UT.g1_i_a4_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNIRM5C62_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__14491\,
            in1 => \N__16015\,
            in2 => \N__14485\,
            in3 => \N__16681\,
            lcout => OPEN,
            ltout => \Lab_UT.g0_3_a3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_3_0_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__14474\,
            in1 => \N__16378\,
            in2 => \N__14449\,
            in3 => \N__14551\,
            lcout => \Lab_UT.g0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIQB3N9_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__18749\,
            in1 => \N__14587\,
            in2 => \N__18600\,
            in3 => \N__23052\,
            lcout => \Lab_UT.N_182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_12_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101010"
        )
    port map (
            in0 => \N__17494\,
            in1 => \N__18562\,
            in2 => \N__23089\,
            in3 => \N__18751\,
            lcout => \Lab_UT.scctrl.g0_1_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIQB3N9_0_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__18750\,
            in1 => \N__14566\,
            in2 => \N__18601\,
            in3 => \N__23053\,
            lcout => \Lab_UT.scctrl.N_182_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g1_i_a4_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__21478\,
            in1 => \N__21529\,
            in2 => \N__17610\,
            in3 => \N__14537\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.a2b.N_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_3_a3_0_3_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__14713\,
            in1 => \N__14560\,
            in2 => \N__14554\,
            in3 => \N__17882\,
            lcout => \Lab_UT.scdp.a2b.g0_3_a3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIESKOU_3_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__21477\,
            in1 => \N__21528\,
            in2 => \_gnd_net_\,
            in3 => \N__14536\,
            lcout => \Lab_UT.scctrl.next_state_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_a13_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19560\,
            in1 => \N__23051\,
            in2 => \N__16230\,
            in3 => \N__19090\,
            lcout => \Lab_UT.scdp.a2b.N_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIOBJ7V_3_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__21479\,
            in1 => \N__21530\,
            in2 => \N__20282\,
            in3 => \N__14538\,
            lcout => \Lab_UT.scctrl.next_state_rst_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_3_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011111010"
        )
    port map (
            in0 => \N__18325\,
            in1 => \N__16675\,
            in2 => \N__20093\,
            in3 => \N__14611\,
            lcout => \Lab_UT.scctrl.N_6_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNI3PVB9_2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20530\,
            in1 => \N__18543\,
            in2 => \N__19553\,
            in3 => \N__18720\,
            lcout => \Lab_UT.state_2_RNI3PVB9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_14_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111111"
        )
    port map (
            in0 => \N__18719\,
            in1 => \N__19180\,
            in2 => \N__18589\,
            in3 => \N__21714\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_9_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__19679\,
            in1 => \_gnd_net_\,
            in2 => \N__14614\,
            in3 => \N__17476\,
            lcout => \Lab_UT.scctrl.g0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_3_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__18982\,
            in1 => \N__14605\,
            in2 => \N__15013\,
            in3 => \N__14596\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_i_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_1_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001110"
        )
    port map (
            in0 => \N__20052\,
            in1 => \N__20341\,
            in2 => \N__14590\,
            in3 => \N__18236\,
            lcout => \Lab_UT.scctrl.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNI1IP99_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__18721\,
            in1 => \N__19678\,
            in2 => \N__18590\,
            in3 => \N__21715\,
            lcout => \Lab_UT.scctrl.N_8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNI5GLD_3_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20487\,
            in2 => \_gnd_net_\,
            in3 => \N__17475\,
            lcout => \Lab_UT.scctrl.un6_sccDecrypt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNI67CB7_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__21408\,
            in1 => \N__23062\,
            in2 => \_gnd_net_\,
            in3 => \N__19096\,
            lcout => \Lab_UT.scctrl.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep2_RNIP9684_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001111"
        )
    port map (
            in0 => \N__22253\,
            in1 => \N__20537\,
            in2 => \N__22102\,
            in3 => \N__18729\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep2_RNIRU4BD_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100011111100"
        )
    port map (
            in0 => \N__16581\,
            in1 => \N__18572\,
            in2 => \N__14578\,
            in3 => \N__20990\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_RNIL9QO21_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16693\,
            in1 => \N__14575\,
            in2 => \N__14569\,
            in3 => \N__17897\,
            lcout => \Lab_UT.scctrl.next_state_rst_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_RNIJN409_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__18728\,
            in1 => \N__20531\,
            in2 => \N__22304\,
            in3 => \N__18571\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_1_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep2_RNIEANJ9_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__17575\,
            in1 => \N__22096\,
            in2 => \N__14716\,
            in3 => \N__21189\,
            lcout => \Lab_UT.next_state_rst_1_3\,
            ltout => \Lab_UT.next_state_rst_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNO_0_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101001111"
        )
    port map (
            in0 => \N__21409\,
            in1 => \N__23063\,
            in2 => \N__14704\,
            in3 => \N__19097\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_0_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__20991\,
            in1 => \N__14700\,
            in2 => \N__14680\,
            in3 => \N__17898\,
            lcout => \Lab_UT.scctrl.next_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22648\,
            ce => \N__14791\,
            sr => \N__18084\
        );

    \Lab_UT.scctrl.state_ret_14_RNITPFM7_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011111"
        )
    port map (
            in0 => \N__23078\,
            in1 => \N__21397\,
            in2 => \N__21735\,
            in3 => \N__19101\,
            lcout => \Lab_UT.next_state_rst_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNIRVOO_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21398\,
            in1 => \N__21668\,
            in2 => \_gnd_net_\,
            in3 => \N__23079\,
            lcout => led_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111110001"
        )
    port map (
            in0 => \N__17218\,
            in1 => \N__14641\,
            in2 => \N__17119\,
            in3 => \N__17182\,
            lcout => \Lab_UT.scctrl.next_state_rst_0_3_N_6_1\,
            ltout => \Lab_UT.scctrl.next_state_rst_0_3_N_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_5_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011111"
        )
    port map (
            in0 => \N__20363\,
            in1 => \_gnd_net_\,
            in2 => \N__14629\,
            in3 => \N__14814\,
            lcout => \Lab_UT.scctrl.g0_i_m4_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_RNIOJNB3_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__21196\,
            in1 => \N__21942\,
            in2 => \N__14752\,
            in3 => \N__21021\,
            lcout => \Lab_UT.scctrl.g0_i_2_0\,
            ltout => \Lab_UT.scctrl.g0_i_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_RNI3MOQ41_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__20364\,
            in1 => \N__14805\,
            in2 => \N__14626\,
            in3 => \N__17708\,
            lcout => \Lab_UT.scctrl.next_state_rst_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__17709\,
            in1 => \N__20365\,
            in2 => \N__14818\,
            in3 => \N__14806\,
            lcout => next_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22642\,
            ce => \N__14794\,
            sr => \N__18086\
        );

    \Lab_UT.scctrl.state_ret_14_RNI4BIC_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21399\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21669\,
            lcout => \Lab_UT.scctrl.g0_i_a8_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep1_RNI2D76_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19834\,
            in2 => \_gnd_net_\,
            in3 => \N__19219\,
            lcout => \Lab_UT.scctrl.G_21_i_a7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_2_3_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__17446\,
            in1 => \N__19107\,
            in2 => \N__23095\,
            in3 => \N__21022\,
            lcout => \Lab_UT.scctrl.N_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_1_3_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__21688\,
            in1 => \N__18626\,
            in2 => \N__22801\,
            in3 => \N__18748\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_0_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__19666\,
            in1 => \N__14743\,
            in2 => \N__14737\,
            in3 => \N__17442\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_1_0_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_3_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__18326\,
            in1 => \N__20284\,
            in2 => \N__14734\,
            in3 => \N__19835\,
            lcout => \Lab_UT.scctrl.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22636\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNI8TAR_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20488\,
            in1 => \N__23086\,
            in2 => \N__19691\,
            in3 => \N__17441\,
            lcout => \Lab_UT.scctrl.next_state75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20631\,
            lcout => \Lab_UT.state_i_3_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22636\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_3_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001010001010"
        )
    port map (
            in0 => \N__17731\,
            in1 => \N__19963\,
            in2 => \N__18332\,
            in3 => \N__17926\,
            lcout => \Lab_UT.scctrl.N_223_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22631\,
            ce => 'H',
            sr => \N__18057\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_9_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19961\,
            in1 => \N__18315\,
            in2 => \_gnd_net_\,
            in3 => \N__17367\,
            lcout => \Lab_UT.scctrl.N_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNO_3_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18952\,
            in2 => \N__18331\,
            in3 => \N__19962\,
            lcout => \Lab_UT.scctrl.N_12_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_3_RNI95RN_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21769\,
            in1 => \N__23087\,
            in2 => \_gnd_net_\,
            in3 => \N__15001\,
            lcout => \Lab_UT.scctrl.next_state73\,
            ltout => \Lab_UT.scctrl.next_state73_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_3_RNII68F41_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14908\,
            in2 => \N__14989\,
            in3 => \N__14981\,
            lcout => \Lab_UT.state_ret_3_RNII68F41_0\,
            ltout => \Lab_UT.state_ret_3_RNII68F41_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.k2l.q_0_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__15223\,
            in1 => \N__14943\,
            in2 => \N__14950\,
            in3 => \N__15511\,
            lcout => \Lab_UT.scdp.key2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22631\,
            ce => 'H',
            sr => \N__18057\
        );

    \Lab_UT.scdp.k2l.q_1_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__14928\,
            in1 => \N__15224\,
            in2 => \N__15390\,
            in3 => \N__14910\,
            lcout => \Lab_UT.scdp.key2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22631\,
            ce => 'H',
            sr => \N__18057\
        );

    \Lab_UT.scdp.k2l.q_2_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14909\,
            in1 => \N__14886\,
            in2 => \N__15273\,
            in3 => \N__15561\,
            lcout => \Lab_UT.scdp.key2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22631\,
            ce => 'H',
            sr => \N__18057\
        );

    \Lab_UT.scdp.rxdataD.q_1_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010111101111"
        )
    port map (
            in0 => \N__15819\,
            in1 => \N__15705\,
            in2 => \N__15789\,
            in3 => \N__14872\,
            lcout => \Lab_UT.scdp.binValD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22627\,
            ce => 'H',
            sr => \N__18059\
        );

    \Lab_UT.scdp.k0h.q_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__15834\,
            in1 => \N__15364\,
            in2 => \N__15279\,
            in3 => \N__15430\,
            lcout => \Lab_UT.scdp.key0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22627\,
            ce => 'H',
            sr => \N__18059\
        );

    \Lab_UT.scdp.rxdataD.q_2_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010000"
        )
    port map (
            in0 => \N__15820\,
            in1 => \_gnd_net_\,
            in2 => \N__15790\,
            in3 => \N__15706\,
            lcout => \Lab_UT.scdp.binValD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22627\,
            ce => 'H',
            sr => \N__18059\
        );

    \Lab_UT.scdp.k0h.q_2_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__15556\,
            in1 => \N__15528\,
            in2 => \N__15280\,
            in3 => \N__15431\,
            lcout => \Lab_UT.scdp.key0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22627\,
            ce => 'H',
            sr => \N__18059\
        );

    \Lab_UT.scdp.k0h.q_0_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__15510\,
            in1 => \N__15447\,
            in2 => \N__15278\,
            in3 => \N__15429\,
            lcout => \Lab_UT.scdp.key0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22627\,
            ce => 'H',
            sr => \N__18059\
        );

    \Lab_UT.scdp.k0h.q_3_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__15432\,
            in1 => \N__15324\,
            in2 => \N__15411\,
            in3 => \N__15265\,
            lcout => \Lab_UT.scdp.key0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22627\,
            ce => 'H',
            sr => \N__18059\
        );

    \Lab_UT.scdp.k0l.q_1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__15339\,
            in1 => \N__15365\,
            in2 => \N__15281\,
            in3 => \N__15077\,
            lcout => \Lab_UT.scdp.key0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22627\,
            ce => 'H',
            sr => \N__18059\
        );

    \Lab_UT.scdp.k0l.q_3_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__15048\,
            in1 => \N__15325\,
            in2 => \N__15282\,
            in3 => \N__15082\,
            lcout => \Lab_UT.scdp.key0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22623\,
            ce => 'H',
            sr => \N__18061\
        );

    \Lab_UT.scctrl.state_ret_13_RNIH6LF_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21947\,
            in1 => \N__20538\,
            in2 => \N__19704\,
            in3 => \N__17498\,
            lcout => \Lab_UT.scctrl.next_state74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.state_ret_5_rep1_RNIP4DD_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__20059\,
            in1 => \N__18938\,
            in2 => \N__17695\,
            in3 => \N__17359\,
            lcout => \G_23_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIR2DQ_3_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__20454\,
            in1 => \N__23092\,
            in2 => \N__20094\,
            in3 => \N__17501\,
            lcout => \Lab_UT.scctrl.N_12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNIOTIG_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__15984\,
            in1 => \N__19703\,
            in2 => \_gnd_net_\,
            in3 => \N__23093\,
            lcout => \Lab_UT.scctrl.g0_0_i_a8_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_RNI493D_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21445\,
            in1 => \N__21870\,
            in2 => \_gnd_net_\,
            in3 => \N__21783\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_0_i_a8_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_RNIMMAAB_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__15973\,
            in1 => \N__16024\,
            in2 => \N__15964\,
            in3 => \N__21024\,
            lcout => \Lab_UT.scctrl.g0_0_i_3_0\,
            ltout => \Lab_UT.scctrl.g0_0_i_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__15923\,
            in1 => \N__15891\,
            in2 => \N__15961\,
            in3 => \N__15944\,
            lcout => \Lab_UT.state_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_4_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15958\,
            in1 => \N__16048\,
            in2 => \N__18954\,
            in3 => \N__15952\,
            lcout => \Lab_UT.scctrl.g0_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep2_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__15858\,
            in1 => \N__15895\,
            in2 => \N__15928\,
            in3 => \N__15946\,
            lcout => \Lab_UT.scctrl.state_i_3_0_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep1_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__15945\,
            in1 => \N__15924\,
            in2 => \N__15898\,
            in3 => \N__15857\,
            lcout => \Lab_UT.state_i_3_0_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ufifo.tx_fsm.cstate_RNO_0_1_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20806\,
            in1 => \N__16207\,
            in2 => \N__16192\,
            in3 => \N__16170\,
            lcout => \ufifo.tx_fsm.N_60_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep1_RNIR7JL_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22378\,
            in2 => \_gnd_net_\,
            in3 => \N__19292\,
            lcout => \Lab_UT.scctrl.N_127_i_i_a6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20632\,
            lcout => \Lab_UT.state_i_3_2_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_7_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19165\,
            in1 => \N__21388\,
            in2 => \N__23075\,
            in3 => \N__19970\,
            lcout => \Lab_UT.scctrl.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_RNIOI524_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000100010"
        )
    port map (
            in0 => \N__16042\,
            in1 => \N__22319\,
            in2 => \N__16036\,
            in3 => \N__20805\,
            lcout => \Lab_UT.scctrl.N_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNI73HE7_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011101"
        )
    port map (
            in0 => \N__17363\,
            in1 => \N__23022\,
            in2 => \N__21425\,
            in3 => \N__19164\,
            lcout => \Lab_UT.scctrl.g0_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNIP81E9_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__21788\,
            in1 => \N__18624\,
            in2 => \N__22420\,
            in3 => \N__18783\,
            lcout => \Lab_UT.N_5\,
            ltout => \Lab_UT.N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_5_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18367\,
            in2 => \N__16018\,
            in3 => \N__19161\,
            lcout => \Lab_UT.g0_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNIFT4T_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__20061\,
            in1 => \N__19697\,
            in2 => \N__17506\,
            in3 => \N__20229\,
            lcout => \Lab_UT.scctrl.g0_14_mb_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNIDM3F1_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__19538\,
            in1 => \N__22994\,
            in2 => \N__22069\,
            in3 => \N__22402\,
            lcout => \Lab_UT.scctrl.g0_0_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNI5UIN_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__20050\,
            in1 => \N__22407\,
            in2 => \N__22092\,
            in3 => \N__22259\,
            lcout => \Lab_UT.scctrl.N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_8_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__19705\,
            in1 => \N__16393\,
            in2 => \N__16231\,
            in3 => \N__17524\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.a2b.g0_iZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_3_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16387\,
            in1 => \N__16615\,
            in2 => \N__16381\,
            in3 => \N__16609\,
            lcout => \Lab_UT.scdp.a2b.g0_3_a3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.g0_i_a5_1_3_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16371\,
            in1 => \N__16970\,
            in2 => \N__16304\,
            in3 => \N__16560\,
            lcout => OPEN,
            ltout => \Lab_UT.g0_i_a5_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_a13_2_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22406\,
            in1 => \N__19309\,
            in2 => \N__16240\,
            in3 => \N__20791\,
            lcout => \Lab_UT.scdp.a2b.N_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNO_7_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100000000"
        )
    port map (
            in0 => \N__20986\,
            in1 => \N__23011\,
            in2 => \N__19167\,
            in3 => \N__17490\,
            lcout => \Lab_UT.scctrl.N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_o13_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22257\,
            in2 => \_gnd_net_\,
            in3 => \N__20539\,
            lcout => \Lab_UT.scdp.a2b.g1_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_4_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__16667\,
            in1 => \N__16213\,
            in2 => \N__20571\,
            in3 => \N__16603\,
            lcout => \Lab_UT.scctrl.g0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNIPVJ8_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__22416\,
            in1 => \N__22258\,
            in2 => \_gnd_net_\,
            in3 => \N__20540\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_127_i_i_o6_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNI9IKA21_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__17224\,
            in1 => \N__16624\,
            in2 => \N__16684\,
            in3 => \N__16605\,
            lcout => \Lab_UT.scctrl.N_127_i_i_a6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_8_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__17489\,
            in1 => \N__19151\,
            in2 => \N__23072\,
            in3 => \N__20985\,
            lcout => \Lab_UT.scctrl.N_190_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_9_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__16668\,
            in1 => \N__16642\,
            in2 => \N__16636\,
            in3 => \N__16623\,
            lcout => \Lab_UT.scdp.a2b.g0_iZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIDJ6UM_0_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__16604\,
            in1 => \N__16588\,
            in2 => \N__16582\,
            in3 => \N__20984\,
            lcout => \Lab_UT.scctrl.g0_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep1_RNI0TTF2_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__19314\,
            in1 => \N__16561\,
            in2 => \_gnd_net_\,
            in3 => \N__20758\,
            lcout => \Lab_UT.scctrl.next_state_1_i_o2_0_d_1\,
            ltout => \Lab_UT.scctrl.next_state_1_i_o2_0_d_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110011"
        )
    port map (
            in0 => \N__17170\,
            in1 => \N__17148\,
            in2 => \N__16513\,
            in3 => \N__17215\,
            lcout => \Lab_UT.state_ret_8_rep1_RNIJDTUE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_rst_0_3_N_5L8_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16966\,
            in2 => \_gnd_net_\,
            in3 => \N__17076\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_0_3_N_5L8Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep1_RNIKN433_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__19315\,
            in1 => \N__16509\,
            in2 => \N__16450\,
            in3 => \N__16446\,
            lcout => \Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433\,
            ltout => \Lab_UT.scctrl.state_ret_8_rep1_RNIKNZ0Z433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__17149\,
            in1 => \N__17239\,
            in2 => \N__17227\,
            in3 => \N__17110\,
            lcout => \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_7_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000111011"
        )
    port map (
            in0 => \N__17111\,
            in1 => \N__17150\,
            in2 => \N__17178\,
            in3 => \N__17216\,
            lcout => \Lab_UT.scctrl.next_state_rst_0_3_N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUE_2_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__17217\,
            in1 => \N__17174\,
            in2 => \N__17155\,
            in3 => \N__17112\,
            lcout => \Lab_UT.scctrl.state_ret_8_rep1_RNIJDTUEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dk.shifter_ret_2_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__17077\,
            in1 => \_gnd_net_\,
            in2 => \N__16972\,
            in3 => \_gnd_net_\,
            lcout => \resetGen_escKey_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22660\,
            ce => \N__16759\,
            sr => \N__18085\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_6_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110000"
        )
    port map (
            in0 => \N__21191\,
            in1 => \N__22435\,
            in2 => \N__17624\,
            in3 => \N__21015\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_2_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__16729\,
            in1 => \N__16711\,
            in2 => \N__16705\,
            in3 => \N__16702\,
            lcout => \Lab_UT.scctrl.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIBABG4_2_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__20569\,
            in1 => \N__17496\,
            in2 => \N__19554\,
            in3 => \N__18780\,
            lcout => \Lab_UT.scctrl.g0_i_a8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_8_RNI3O64_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__21190\,
            in1 => \N__17625\,
            in2 => \_gnd_net_\,
            in3 => \N__21922\,
            lcout => \Lab_UT.scctrl.g0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNITPFM7_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010111"
        )
    port map (
            in0 => \N__21756\,
            in1 => \N__23091\,
            in2 => \N__21444\,
            in3 => \N__19157\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_rst_0_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNIB361N_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__17611\,
            in1 => \N__17520\,
            in2 => \N__17509\,
            in3 => \N__18175\,
            lcout => \Lab_UT.scctrl.g0_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNIT01T_3_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__17495\,
            in1 => \N__23090\,
            in2 => \N__17368\,
            in3 => \N__20570\,
            lcout => \Lab_UT.scctrl.g0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_2_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__18327\,
            in1 => \N__19877\,
            in2 => \_gnd_net_\,
            in3 => \N__18246\,
            lcout => \Lab_UT.scctrl.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNINBNBI_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__17752\,
            in1 => \N__17299\,
            in2 => \N__17293\,
            in3 => \N__18625\,
            lcout => \Lab_UT.scctrl.g0_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNITQ09E1_1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100110011"
        )
    port map (
            in0 => \N__17284\,
            in1 => \N__17681\,
            in2 => \N__17275\,
            in3 => \N__19876\,
            lcout => \Lab_UT.scctrl.g2\,
            ltout => \Lab_UT.scctrl.g2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIM7FBH2_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010110000"
        )
    port map (
            in0 => \N__19878\,
            in1 => \N__18422\,
            in2 => \N__17266\,
            in3 => \N__18102\,
            lcout => \Lab_UT.scctrl.N_223_1_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__19880\,
            in1 => \N__17263\,
            in2 => \N__17691\,
            in3 => \N__17257\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_222i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101111"
        )
    port map (
            in0 => \N__18922\,
            in1 => \N__17908\,
            in2 => \N__17248\,
            in3 => \N__17245\,
            lcout => \Lab_UT_scctrl_N_221_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIDKJEO1_3_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010001100"
        )
    port map (
            in0 => \N__19879\,
            in1 => \N__17730\,
            in2 => \N__18336\,
            in3 => \N__17925\,
            lcout => \Lab_UT.scctrl.N_223_2_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100111"
        )
    port map (
            in0 => \N__19967\,
            in1 => \N__17902\,
            in2 => \N__18443\,
            in3 => \N__17863\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_i_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__17632\,
            in1 => \N__17851\,
            in2 => \N__17845\,
            in3 => \N__17716\,
            lcout => led_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNITPFM7_1_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__19149\,
            in1 => \N__21432\,
            in2 => \N__21792\,
            in3 => \N__23074\,
            lcout => \Lab_UT.scctrl.N_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIEUO38_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110001101"
        )
    port map (
            in0 => \N__19875\,
            in1 => \N__18346\,
            in2 => \N__20349\,
            in3 => \N__19148\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_18_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNIE2CTO_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000111"
        )
    port map (
            in0 => \N__19964\,
            in1 => \N__17743\,
            in2 => \N__17734\,
            in3 => \N__18802\,
            lcout => \Lab_UT.scctrl.next_stateZ0Z_2\,
            ltout => \Lab_UT.scctrl.next_stateZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20267\,
            in2 => \N__17719\,
            in3 => \N__19966\,
            lcout => \Lab_UT.scctrl.N_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_15_RNO_3_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110101111"
        )
    port map (
            in0 => \N__19965\,
            in1 => \N__17710\,
            in2 => \N__17685\,
            in3 => \N__17638\,
            lcout => \Lab_UT.scctrl.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNI6VDS_0_2_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__19552\,
            in1 => \N__20574\,
            in2 => \N__22191\,
            in3 => \N__23077\,
            lcout => \Lab_UT.scctrl.g1_i_a7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_RNO_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000111"
        )
    port map (
            in0 => \N__20268\,
            in1 => \N__19968\,
            in2 => \N__18337\,
            in3 => \N__18247\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.next_state_i_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18223\,
            in3 => \N__18951\,
            lcout => \Lab_UT.state_i_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNI6VDS_2_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19551\,
            in1 => \N__20572\,
            in2 => \N__22190\,
            in3 => \N__23076\,
            lcout => \Lab_UT.scctrl.next_state71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIR2DQ_2_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19530\,
            in1 => \N__21943\,
            in2 => \N__22192\,
            in3 => \N__21770\,
            lcout => \Lab_UT.scctrl.next_state72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNIPVJ8_0_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__22415\,
            in1 => \N__22152\,
            in2 => \_gnd_net_\,
            in3 => \N__20573\,
            lcout => \Lab_UT.scctrl.g4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.EmsBitsSl_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18140\,
            lcout => \Lab_UT.sccEmsBitsSl\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22632\,
            ce => 'H',
            sr => \N__18062\
        );

    \Lab_UT.scctrl.state_ret_6_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000001010001010"
        )
    port map (
            in0 => \N__18118\,
            in1 => \N__19969\,
            in2 => \N__18450\,
            in3 => \N__18109\,
            lcout => \Lab_UT.scctrl.N_223_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22632\,
            ce => 'H',
            sr => \N__18062\
        );

    \Lab_UT.scctrl.state_1_RNO_5_0_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__21928\,
            in1 => \N__20565\,
            in2 => \N__22332\,
            in3 => \N__18784\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_0_i_a8_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_1_0_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__18379\,
            in1 => \N__18373\,
            in2 => \N__18472\,
            in3 => \N__18628\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_38_0_a3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_0_0_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__21562\,
            in1 => \N__18469\,
            in2 => \N__18454\,
            in3 => \N__21020\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_38_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_0_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__18451\,
            in1 => \N__18869\,
            in2 => \N__18382\,
            in3 => \N__20070\,
            lcout => \Lab_UT.state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_6_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__21929\,
            in1 => \N__21185\,
            in2 => \_gnd_net_\,
            in3 => \N__21019\,
            lcout => \Lab_UT.scctrl.N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_4_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100101111"
        )
    port map (
            in0 => \N__22920\,
            in1 => \N__21407\,
            in2 => \N__20257\,
            in3 => \N__19156\,
            lcout => \Lab_UT.scctrl.g0_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_a9_1_0_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__19521\,
            in1 => \N__20564\,
            in2 => \N__22331\,
            in3 => \N__22919\,
            lcout => \Lab_UT.scdp.a2b.g0_i_a9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_9_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20556\,
            in1 => \N__19658\,
            in2 => \N__23019\,
            in3 => \N__22326\,
            lcout => \Lab_UT.scctrl.g0_0_i_a8_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__21975\,
            in1 => \N__18858\,
            in2 => \_gnd_net_\,
            in3 => \N__20019\,
            lcout => OPEN,
            ltout => \Lab_UT.scdp.a2b.g0_iZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scdp.a2b.g0_i_2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__19319\,
            in1 => \N__22324\,
            in2 => \N__18358\,
            in3 => \N__19243\,
            lcout => \Lab_UT.scdp.a2b.g0_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_15_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__22323\,
            in1 => \N__20020\,
            in2 => \N__19323\,
            in3 => \N__20555\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_7_a13_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_12_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18620\,
            in2 => \N__18973\,
            in3 => \N__18773\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_5_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19371\,
            in1 => \N__19342\,
            in2 => \N__18970\,
            in3 => \N__18790\,
            lcout => \Lab_UT.scctrl.g0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_11_RNI7NLQ7_0_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__20554\,
            in1 => \N__22325\,
            in2 => \N__19393\,
            in3 => \N__19168\,
            lcout => \Lab_UT.scctrl.N_9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_0_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22788\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNIFKMJ3_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22421\,
            in1 => \N__18814\,
            in2 => \N__20815\,
            in3 => \N__22073\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_10_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNI0K8F7_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__21961\,
            in1 => \N__21175\,
            in2 => \N__18805\,
            in3 => \N__20982\,
            lcout => \Lab_UT.scctrl.g1_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_13_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__19996\,
            in1 => \N__21174\,
            in2 => \N__22094\,
            in3 => \N__20981\,
            lcout => \Lab_UT.scctrl.N_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_0_RNIN6IE9_1_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__21787\,
            in1 => \N__18765\,
            in2 => \N__18643\,
            in3 => \N__18616\,
            lcout => \Lab_UT.scctrl.N_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNIBRA17_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__19997\,
            in1 => \N__19429\,
            in2 => \N__21207\,
            in3 => \N__20983\,
            lcout => \Lab_UT.scctrl.G_21_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNO_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__19379\,
            in1 => \N__20270\,
            in2 => \_gnd_net_\,
            in3 => \N__19344\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_24_i_a4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__19408\,
            in1 => \N__21454\,
            in2 => \N__19396\,
            in3 => \N__20641\,
            lcout => \Lab_UT.N_169_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19381\,
            in1 => \N__19717\,
            in2 => \N__19360\,
            in3 => \N__19345\,
            lcout => \Lab_UT.state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_2_RNIGC1Q_0_2_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22955\,
            in1 => \N__19992\,
            in2 => \_gnd_net_\,
            in3 => \N__19486\,
            lcout => \Lab_UT.scctrl.G_21_i_a7_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_9_RNIPD53P_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19380\,
            in1 => \N__19716\,
            in2 => \N__19359\,
            in3 => \N__19343\,
            lcout => \Lab_UT.scctrl.N_4ctr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.nibbleIn1_RNO_16_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__22956\,
            in1 => \N__19487\,
            in2 => \N__19327\,
            in3 => \N__19239\,
            lcout => \Lab_UT.scctrl.g0_1_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_15_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__19485\,
            in1 => \_gnd_net_\,
            in2 => \N__20069\,
            in3 => \N__22957\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.g0_i_a7_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_10_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__22301\,
            in1 => \N__20578\,
            in2 => \N__19171\,
            in3 => \N__19155\,
            lcout => \Lab_UT.scctrl.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNO_4_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21206\,
            in2 => \_gnd_net_\,
            in3 => \N__21025\,
            lcout => \Lab_UT.scctrl.N_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNO_8_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19621\,
            in2 => \_gnd_net_\,
            in3 => \N__21948\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.G_24_i_o3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNO_5_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111010"
        )
    port map (
            in0 => \N__22297\,
            in1 => \N__20830\,
            in2 => \N__20818\,
            in3 => \N__20814\,
            lcout => OPEN,
            ltout => \Lab_UT.scctrl.N_6_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNO_1_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19972\,
            in1 => \N__20350\,
            in2 => \N__20650\,
            in3 => \N__20647\,
            lcout => \Lab_UT.scctrl.N_8_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20611\,
            lcout => \Lab_UT.state_i_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNIQT9P_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__19971\,
            in1 => \N__21290\,
            in2 => \N__21793\,
            in3 => \N__23002\,
            lcout => \Lab_UT.scctrl.G_23_0_a9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_RNI19C4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22296\,
            in1 => \N__19628\,
            in2 => \_gnd_net_\,
            in3 => \N__20575\,
            lcout => \Lab_UT.scctrl.g0_i_a8_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.next_state_RNIGKIO_2_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__20348\,
            in1 => \N__20269\,
            in2 => \_gnd_net_\,
            in3 => \N__19998\,
            lcout => \Lab_UT.scctrl.G_21_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_3_3_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__19654\,
            in1 => \N__21951\,
            in2 => \N__19550\,
            in3 => \N__23018\,
            lcout => \Lab_UT.scctrl.g0_i_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.state_ret_5_fast_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22789\,
            lcout => rst_i_3_fast,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_7_RNO_13_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__21362\,
            in1 => \N__22077\,
            in2 => \_gnd_net_\,
            in3 => \N__21789\,
            lcout => \Lab_UT.scctrl.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_13_rep2_RNITKTS_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__22423\,
            in1 => \N__22327\,
            in2 => \N__22095\,
            in3 => \N__21976\,
            lcout => \Lab_UT.scctrl.g1_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_1_RNO_3_0_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__21363\,
            in1 => \N__21923\,
            in2 => \N__21802\,
            in3 => \N__21790\,
            lcout => \Lab_UT.scctrl.state_1_RNO_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_14_RNO_2_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__21556\,
            in1 => \N__21547\,
            in2 => \N__21508\,
            in3 => \N__21490\,
            lcout => \Lab_UT.scctrl.N_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.scctrl.state_ret_6_RNIBMV1_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21324\,
            in2 => \_gnd_net_\,
            in3 => \N__21253\,
            lcout => led_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
