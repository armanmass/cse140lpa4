// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Jun 3 2019 04:43:08

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__23809;
    wire N__23808;
    wire N__23807;
    wire N__23800;
    wire N__23799;
    wire N__23798;
    wire N__23791;
    wire N__23790;
    wire N__23789;
    wire N__23782;
    wire N__23781;
    wire N__23780;
    wire N__23773;
    wire N__23772;
    wire N__23771;
    wire N__23764;
    wire N__23763;
    wire N__23762;
    wire N__23755;
    wire N__23754;
    wire N__23753;
    wire N__23746;
    wire N__23745;
    wire N__23744;
    wire N__23737;
    wire N__23736;
    wire N__23735;
    wire N__23728;
    wire N__23727;
    wire N__23726;
    wire N__23709;
    wire N__23708;
    wire N__23707;
    wire N__23706;
    wire N__23705;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23697;
    wire N__23696;
    wire N__23695;
    wire N__23692;
    wire N__23691;
    wire N__23690;
    wire N__23687;
    wire N__23676;
    wire N__23673;
    wire N__23672;
    wire N__23669;
    wire N__23668;
    wire N__23663;
    wire N__23660;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23638;
    wire N__23635;
    wire N__23630;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23614;
    wire N__23607;
    wire N__23606;
    wire N__23605;
    wire N__23604;
    wire N__23601;
    wire N__23600;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23589;
    wire N__23586;
    wire N__23581;
    wire N__23574;
    wire N__23573;
    wire N__23572;
    wire N__23569;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23525;
    wire N__23524;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23513;
    wire N__23510;
    wire N__23509;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23505;
    wire N__23504;
    wire N__23503;
    wire N__23502;
    wire N__23501;
    wire N__23500;
    wire N__23499;
    wire N__23498;
    wire N__23497;
    wire N__23496;
    wire N__23495;
    wire N__23494;
    wire N__23493;
    wire N__23492;
    wire N__23491;
    wire N__23490;
    wire N__23489;
    wire N__23488;
    wire N__23487;
    wire N__23484;
    wire N__23481;
    wire N__23478;
    wire N__23475;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23463;
    wire N__23458;
    wire N__23455;
    wire N__23454;
    wire N__23453;
    wire N__23452;
    wire N__23449;
    wire N__23448;
    wire N__23445;
    wire N__23444;
    wire N__23443;
    wire N__23442;
    wire N__23441;
    wire N__23440;
    wire N__23439;
    wire N__23438;
    wire N__23435;
    wire N__23434;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23426;
    wire N__23425;
    wire N__23422;
    wire N__23421;
    wire N__23416;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23394;
    wire N__23393;
    wire N__23392;
    wire N__23391;
    wire N__23390;
    wire N__23389;
    wire N__23388;
    wire N__23381;
    wire N__23378;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23352;
    wire N__23351;
    wire N__23350;
    wire N__23349;
    wire N__23348;
    wire N__23345;
    wire N__23334;
    wire N__23323;
    wire N__23318;
    wire N__23305;
    wire N__23298;
    wire N__23293;
    wire N__23280;
    wire N__23273;
    wire N__23264;
    wire N__23261;
    wire N__23252;
    wire N__23247;
    wire N__23242;
    wire N__23239;
    wire N__23230;
    wire N__23211;
    wire N__23210;
    wire N__23209;
    wire N__23208;
    wire N__23203;
    wire N__23202;
    wire N__23199;
    wire N__23198;
    wire N__23197;
    wire N__23196;
    wire N__23195;
    wire N__23192;
    wire N__23191;
    wire N__23190;
    wire N__23189;
    wire N__23188;
    wire N__23187;
    wire N__23186;
    wire N__23185;
    wire N__23184;
    wire N__23183;
    wire N__23182;
    wire N__23181;
    wire N__23180;
    wire N__23179;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23162;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23150;
    wire N__23149;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23129;
    wire N__23128;
    wire N__23127;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23119;
    wire N__23118;
    wire N__23117;
    wire N__23112;
    wire N__23109;
    wire N__23108;
    wire N__23105;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23044;
    wire N__23039;
    wire N__23036;
    wire N__23023;
    wire N__23010;
    wire N__23005;
    wire N__23000;
    wire N__22993;
    wire N__22980;
    wire N__22977;
    wire N__22976;
    wire N__22975;
    wire N__22972;
    wire N__22971;
    wire N__22970;
    wire N__22969;
    wire N__22968;
    wire N__22967;
    wire N__22966;
    wire N__22965;
    wire N__22964;
    wire N__22963;
    wire N__22962;
    wire N__22961;
    wire N__22958;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22944;
    wire N__22941;
    wire N__22934;
    wire N__22927;
    wire N__22922;
    wire N__22919;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22877;
    wire N__22872;
    wire N__22865;
    wire N__22860;
    wire N__22857;
    wire N__22842;
    wire N__22841;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22829;
    wire N__22828;
    wire N__22827;
    wire N__22826;
    wire N__22825;
    wire N__22824;
    wire N__22823;
    wire N__22822;
    wire N__22821;
    wire N__22820;
    wire N__22819;
    wire N__22816;
    wire N__22815;
    wire N__22808;
    wire N__22805;
    wire N__22804;
    wire N__22803;
    wire N__22802;
    wire N__22793;
    wire N__22792;
    wire N__22791;
    wire N__22790;
    wire N__22789;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22769;
    wire N__22766;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22747;
    wire N__22742;
    wire N__22741;
    wire N__22738;
    wire N__22737;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22700;
    wire N__22699;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22687;
    wire N__22682;
    wire N__22679;
    wire N__22670;
    wire N__22665;
    wire N__22658;
    wire N__22641;
    wire N__22638;
    wire N__22637;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22585;
    wire N__22584;
    wire N__22583;
    wire N__22582;
    wire N__22581;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22564;
    wire N__22563;
    wire N__22562;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22548;
    wire N__22543;
    wire N__22542;
    wire N__22541;
    wire N__22540;
    wire N__22539;
    wire N__22538;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22485;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22463;
    wire N__22462;
    wire N__22461;
    wire N__22460;
    wire N__22459;
    wire N__22458;
    wire N__22455;
    wire N__22454;
    wire N__22451;
    wire N__22450;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22442;
    wire N__22441;
    wire N__22440;
    wire N__22437;
    wire N__22436;
    wire N__22433;
    wire N__22432;
    wire N__22429;
    wire N__22428;
    wire N__22425;
    wire N__22424;
    wire N__22421;
    wire N__22420;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22359;
    wire N__22356;
    wire N__22351;
    wire N__22342;
    wire N__22339;
    wire N__22334;
    wire N__22331;
    wire N__22326;
    wire N__22323;
    wire N__22316;
    wire N__22313;
    wire N__22308;
    wire N__22303;
    wire N__22296;
    wire N__22293;
    wire N__22292;
    wire N__22291;
    wire N__22290;
    wire N__22289;
    wire N__22288;
    wire N__22287;
    wire N__22286;
    wire N__22285;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22275;
    wire N__22270;
    wire N__22269;
    wire N__22268;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22260;
    wire N__22259;
    wire N__22258;
    wire N__22257;
    wire N__22256;
    wire N__22251;
    wire N__22250;
    wire N__22247;
    wire N__22242;
    wire N__22237;
    wire N__22236;
    wire N__22235;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22210;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22202;
    wire N__22201;
    wire N__22200;
    wire N__22199;
    wire N__22198;
    wire N__22197;
    wire N__22196;
    wire N__22195;
    wire N__22194;
    wire N__22193;
    wire N__22192;
    wire N__22191;
    wire N__22190;
    wire N__22189;
    wire N__22188;
    wire N__22187;
    wire N__22186;
    wire N__22183;
    wire N__22178;
    wire N__22177;
    wire N__22176;
    wire N__22175;
    wire N__22170;
    wire N__22165;
    wire N__22158;
    wire N__22155;
    wire N__22150;
    wire N__22141;
    wire N__22134;
    wire N__22131;
    wire N__22126;
    wire N__22123;
    wire N__22116;
    wire N__22109;
    wire N__22104;
    wire N__22097;
    wire N__22090;
    wire N__22083;
    wire N__22076;
    wire N__22059;
    wire N__22058;
    wire N__22057;
    wire N__22056;
    wire N__22055;
    wire N__22054;
    wire N__22053;
    wire N__22052;
    wire N__22051;
    wire N__22050;
    wire N__22047;
    wire N__22046;
    wire N__22045;
    wire N__22044;
    wire N__22043;
    wire N__22042;
    wire N__22041;
    wire N__22038;
    wire N__22037;
    wire N__22036;
    wire N__22035;
    wire N__22034;
    wire N__22033;
    wire N__22032;
    wire N__22031;
    wire N__22030;
    wire N__22029;
    wire N__22028;
    wire N__22027;
    wire N__22024;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22003;
    wire N__21998;
    wire N__21997;
    wire N__21996;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21990;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21976;
    wire N__21975;
    wire N__21974;
    wire N__21973;
    wire N__21972;
    wire N__21971;
    wire N__21966;
    wire N__21965;
    wire N__21962;
    wire N__21961;
    wire N__21960;
    wire N__21957;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21945;
    wire N__21938;
    wire N__21929;
    wire N__21928;
    wire N__21921;
    wire N__21910;
    wire N__21905;
    wire N__21896;
    wire N__21889;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21875;
    wire N__21874;
    wire N__21873;
    wire N__21872;
    wire N__21867;
    wire N__21864;
    wire N__21859;
    wire N__21858;
    wire N__21855;
    wire N__21854;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21831;
    wire N__21828;
    wire N__21819;
    wire N__21818;
    wire N__21817;
    wire N__21816;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21787;
    wire N__21780;
    wire N__21775;
    wire N__21768;
    wire N__21761;
    wire N__21758;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21728;
    wire N__21725;
    wire N__21724;
    wire N__21723;
    wire N__21722;
    wire N__21721;
    wire N__21718;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21710;
    wire N__21709;
    wire N__21708;
    wire N__21707;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21692;
    wire N__21687;
    wire N__21682;
    wire N__21677;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21653;
    wire N__21650;
    wire N__21645;
    wire N__21640;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21623;
    wire N__21622;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21597;
    wire N__21594;
    wire N__21593;
    wire N__21590;
    wire N__21589;
    wire N__21588;
    wire N__21585;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21570;
    wire N__21567;
    wire N__21562;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21537;
    wire N__21536;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21521;
    wire N__21520;
    wire N__21519;
    wire N__21518;
    wire N__21515;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21503;
    wire N__21502;
    wire N__21501;
    wire N__21500;
    wire N__21499;
    wire N__21498;
    wire N__21497;
    wire N__21496;
    wire N__21495;
    wire N__21492;
    wire N__21489;
    wire N__21484;
    wire N__21481;
    wire N__21480;
    wire N__21479;
    wire N__21472;
    wire N__21467;
    wire N__21464;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21437;
    wire N__21432;
    wire N__21417;
    wire N__21416;
    wire N__21415;
    wire N__21414;
    wire N__21413;
    wire N__21412;
    wire N__21411;
    wire N__21410;
    wire N__21409;
    wire N__21408;
    wire N__21405;
    wire N__21404;
    wire N__21403;
    wire N__21402;
    wire N__21399;
    wire N__21392;
    wire N__21391;
    wire N__21390;
    wire N__21389;
    wire N__21388;
    wire N__21381;
    wire N__21378;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21370;
    wire N__21369;
    wire N__21366;
    wire N__21365;
    wire N__21364;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21342;
    wire N__21339;
    wire N__21334;
    wire N__21333;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21321;
    wire N__21318;
    wire N__21317;
    wire N__21316;
    wire N__21315;
    wire N__21314;
    wire N__21309;
    wire N__21306;
    wire N__21305;
    wire N__21300;
    wire N__21297;
    wire N__21288;
    wire N__21283;
    wire N__21280;
    wire N__21275;
    wire N__21272;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21243;
    wire N__21236;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21188;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21150;
    wire N__21149;
    wire N__21148;
    wire N__21147;
    wire N__21146;
    wire N__21145;
    wire N__21144;
    wire N__21143;
    wire N__21142;
    wire N__21141;
    wire N__21140;
    wire N__21139;
    wire N__21138;
    wire N__21137;
    wire N__21136;
    wire N__21135;
    wire N__21134;
    wire N__21133;
    wire N__21132;
    wire N__21131;
    wire N__21130;
    wire N__21129;
    wire N__21128;
    wire N__21127;
    wire N__21126;
    wire N__21125;
    wire N__21124;
    wire N__21123;
    wire N__21122;
    wire N__21121;
    wire N__21120;
    wire N__21119;
    wire N__21118;
    wire N__21117;
    wire N__21116;
    wire N__21115;
    wire N__21114;
    wire N__21113;
    wire N__21112;
    wire N__21111;
    wire N__21110;
    wire N__21109;
    wire N__21108;
    wire N__21107;
    wire N__21106;
    wire N__21105;
    wire N__21104;
    wire N__21103;
    wire N__21102;
    wire N__21101;
    wire N__21100;
    wire N__21099;
    wire N__21098;
    wire N__21097;
    wire N__21096;
    wire N__21095;
    wire N__21094;
    wire N__21093;
    wire N__21092;
    wire N__21091;
    wire N__21090;
    wire N__21089;
    wire N__21088;
    wire N__21087;
    wire N__21086;
    wire N__21085;
    wire N__21084;
    wire N__21083;
    wire N__21082;
    wire N__21081;
    wire N__21080;
    wire N__21079;
    wire N__21078;
    wire N__21077;
    wire N__21076;
    wire N__21075;
    wire N__21074;
    wire N__21073;
    wire N__21072;
    wire N__21071;
    wire N__21070;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20900;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20869;
    wire N__20862;
    wire N__20859;
    wire N__20858;
    wire N__20857;
    wire N__20856;
    wire N__20855;
    wire N__20854;
    wire N__20853;
    wire N__20852;
    wire N__20851;
    wire N__20850;
    wire N__20849;
    wire N__20848;
    wire N__20847;
    wire N__20846;
    wire N__20845;
    wire N__20844;
    wire N__20843;
    wire N__20842;
    wire N__20841;
    wire N__20840;
    wire N__20839;
    wire N__20838;
    wire N__20837;
    wire N__20836;
    wire N__20835;
    wire N__20834;
    wire N__20833;
    wire N__20832;
    wire N__20831;
    wire N__20830;
    wire N__20829;
    wire N__20828;
    wire N__20827;
    wire N__20826;
    wire N__20825;
    wire N__20824;
    wire N__20823;
    wire N__20822;
    wire N__20821;
    wire N__20820;
    wire N__20819;
    wire N__20818;
    wire N__20817;
    wire N__20816;
    wire N__20815;
    wire N__20814;
    wire N__20813;
    wire N__20812;
    wire N__20811;
    wire N__20810;
    wire N__20809;
    wire N__20808;
    wire N__20807;
    wire N__20804;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20690;
    wire N__20687;
    wire N__20686;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20664;
    wire N__20663;
    wire N__20662;
    wire N__20661;
    wire N__20658;
    wire N__20657;
    wire N__20656;
    wire N__20655;
    wire N__20652;
    wire N__20651;
    wire N__20648;
    wire N__20647;
    wire N__20644;
    wire N__20643;
    wire N__20642;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20609;
    wire N__20606;
    wire N__20605;
    wire N__20596;
    wire N__20591;
    wire N__20586;
    wire N__20585;
    wire N__20578;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20541;
    wire N__20538;
    wire N__20535;
    wire N__20532;
    wire N__20529;
    wire N__20528;
    wire N__20525;
    wire N__20524;
    wire N__20523;
    wire N__20522;
    wire N__20521;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20513;
    wire N__20512;
    wire N__20509;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20491;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20475;
    wire N__20472;
    wire N__20457;
    wire N__20456;
    wire N__20453;
    wire N__20452;
    wire N__20451;
    wire N__20448;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20434;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20419;
    wire N__20414;
    wire N__20411;
    wire N__20404;
    wire N__20399;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20358;
    wire N__20355;
    wire N__20354;
    wire N__20351;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20288;
    wire N__20287;
    wire N__20286;
    wire N__20285;
    wire N__20284;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20269;
    wire N__20268;
    wire N__20267;
    wire N__20262;
    wire N__20259;
    wire N__20258;
    wire N__20253;
    wire N__20252;
    wire N__20251;
    wire N__20250;
    wire N__20247;
    wire N__20236;
    wire N__20233;
    wire N__20228;
    wire N__20225;
    wire N__20218;
    wire N__20209;
    wire N__20204;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20183;
    wire N__20182;
    wire N__20181;
    wire N__20180;
    wire N__20179;
    wire N__20178;
    wire N__20177;
    wire N__20176;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20161;
    wire N__20158;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20141;
    wire N__20140;
    wire N__20139;
    wire N__20136;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20118;
    wire N__20115;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20092;
    wire N__20089;
    wire N__20084;
    wire N__20079;
    wire N__20076;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20054;
    wire N__20053;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20045;
    wire N__20040;
    wire N__20039;
    wire N__20038;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20018;
    wire N__20017;
    wire N__20016;
    wire N__20015;
    wire N__20014;
    wire N__20011;
    wire N__20006;
    wire N__20001;
    wire N__19998;
    wire N__19991;
    wire N__19980;
    wire N__19977;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19946;
    wire N__19945;
    wire N__19944;
    wire N__19943;
    wire N__19942;
    wire N__19941;
    wire N__19936;
    wire N__19935;
    wire N__19934;
    wire N__19931;
    wire N__19930;
    wire N__19927;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19907;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19891;
    wire N__19890;
    wire N__19887;
    wire N__19882;
    wire N__19877;
    wire N__19874;
    wire N__19873;
    wire N__19870;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19847;
    wire N__19836;
    wire N__19833;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19815;
    wire N__19814;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19796;
    wire N__19793;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19730;
    wire N__19729;
    wire N__19728;
    wire N__19727;
    wire N__19726;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19687;
    wire N__19682;
    wire N__19681;
    wire N__19676;
    wire N__19671;
    wire N__19670;
    wire N__19669;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19650;
    wire N__19645;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19607;
    wire N__19604;
    wire N__19603;
    wire N__19600;
    wire N__19599;
    wire N__19598;
    wire N__19597;
    wire N__19596;
    wire N__19591;
    wire N__19588;
    wire N__19581;
    wire N__19578;
    wire N__19577;
    wire N__19574;
    wire N__19573;
    wire N__19572;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19553;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19535;
    wire N__19534;
    wire N__19531;
    wire N__19530;
    wire N__19529;
    wire N__19526;
    wire N__19525;
    wire N__19522;
    wire N__19521;
    wire N__19520;
    wire N__19519;
    wire N__19518;
    wire N__19513;
    wire N__19500;
    wire N__19497;
    wire N__19496;
    wire N__19495;
    wire N__19494;
    wire N__19493;
    wire N__19492;
    wire N__19489;
    wire N__19484;
    wire N__19481;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19444;
    wire N__19441;
    wire N__19434;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19391;
    wire N__19390;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19355;
    wire N__19352;
    wire N__19341;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19333;
    wire N__19332;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19317;
    wire N__19316;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19251;
    wire N__19248;
    wire N__19247;
    wire N__19246;
    wire N__19245;
    wire N__19244;
    wire N__19243;
    wire N__19242;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19222;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19157;
    wire N__19156;
    wire N__19155;
    wire N__19154;
    wire N__19153;
    wire N__19152;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19144;
    wire N__19141;
    wire N__19134;
    wire N__19133;
    wire N__19132;
    wire N__19131;
    wire N__19126;
    wire N__19125;
    wire N__19122;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19104;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19054;
    wire N__19049;
    wire N__19042;
    wire N__19035;
    wire N__19032;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__18999;
    wire N__18996;
    wire N__18993;
    wire N__18990;
    wire N__18987;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18966;
    wire N__18963;
    wire N__18960;
    wire N__18957;
    wire N__18954;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18905;
    wire N__18904;
    wire N__18903;
    wire N__18900;
    wire N__18899;
    wire N__18898;
    wire N__18897;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18887;
    wire N__18884;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18865;
    wire N__18862;
    wire N__18861;
    wire N__18858;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18838;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18813;
    wire N__18812;
    wire N__18809;
    wire N__18808;
    wire N__18805;
    wire N__18804;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18789;
    wire N__18788;
    wire N__18787;
    wire N__18786;
    wire N__18785;
    wire N__18784;
    wire N__18783;
    wire N__18782;
    wire N__18781;
    wire N__18780;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18757;
    wire N__18756;
    wire N__18755;
    wire N__18748;
    wire N__18743;
    wire N__18740;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18689;
    wire N__18688;
    wire N__18687;
    wire N__18686;
    wire N__18685;
    wire N__18684;
    wire N__18683;
    wire N__18682;
    wire N__18681;
    wire N__18680;
    wire N__18679;
    wire N__18678;
    wire N__18677;
    wire N__18676;
    wire N__18675;
    wire N__18674;
    wire N__18671;
    wire N__18670;
    wire N__18669;
    wire N__18668;
    wire N__18667;
    wire N__18666;
    wire N__18665;
    wire N__18664;
    wire N__18661;
    wire N__18660;
    wire N__18659;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18647;
    wire N__18642;
    wire N__18633;
    wire N__18624;
    wire N__18623;
    wire N__18606;
    wire N__18595;
    wire N__18590;
    wire N__18587;
    wire N__18580;
    wire N__18577;
    wire N__18576;
    wire N__18575;
    wire N__18574;
    wire N__18571;
    wire N__18566;
    wire N__18561;
    wire N__18558;
    wire N__18551;
    wire N__18546;
    wire N__18543;
    wire N__18534;
    wire N__18533;
    wire N__18532;
    wire N__18531;
    wire N__18526;
    wire N__18521;
    wire N__18518;
    wire N__18517;
    wire N__18516;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18501;
    wire N__18496;
    wire N__18489;
    wire N__18488;
    wire N__18485;
    wire N__18484;
    wire N__18483;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18468;
    wire N__18459;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18441;
    wire N__18440;
    wire N__18439;
    wire N__18438;
    wire N__18437;
    wire N__18434;
    wire N__18433;
    wire N__18432;
    wire N__18431;
    wire N__18430;
    wire N__18429;
    wire N__18428;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18420;
    wire N__18417;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18406;
    wire N__18399;
    wire N__18396;
    wire N__18395;
    wire N__18392;
    wire N__18387;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18371;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18356;
    wire N__18355;
    wire N__18352;
    wire N__18347;
    wire N__18338;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18315;
    wire N__18312;
    wire N__18307;
    wire N__18304;
    wire N__18301;
    wire N__18296;
    wire N__18291;
    wire N__18282;
    wire N__18279;
    wire N__18278;
    wire N__18277;
    wire N__18276;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18265;
    wire N__18264;
    wire N__18263;
    wire N__18260;
    wire N__18259;
    wire N__18256;
    wire N__18251;
    wire N__18248;
    wire N__18247;
    wire N__18246;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18238;
    wire N__18235;
    wire N__18232;
    wire N__18231;
    wire N__18230;
    wire N__18227;
    wire N__18226;
    wire N__18225;
    wire N__18222;
    wire N__18217;
    wire N__18212;
    wire N__18209;
    wire N__18204;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18182;
    wire N__18177;
    wire N__18174;
    wire N__18169;
    wire N__18166;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18113;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18086;
    wire N__18085;
    wire N__18082;
    wire N__18079;
    wire N__18076;
    wire N__18073;
    wire N__18072;
    wire N__18071;
    wire N__18068;
    wire N__18067;
    wire N__18066;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18058;
    wire N__18055;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18043;
    wire N__18040;
    wire N__18039;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18019;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18004;
    wire N__17999;
    wire N__17994;
    wire N__17991;
    wire N__17988;
    wire N__17983;
    wire N__17976;
    wire N__17973;
    wire N__17968;
    wire N__17955;
    wire N__17952;
    wire N__17951;
    wire N__17950;
    wire N__17949;
    wire N__17948;
    wire N__17945;
    wire N__17936;
    wire N__17931;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17913;
    wire N__17910;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17898;
    wire N__17897;
    wire N__17896;
    wire N__17895;
    wire N__17894;
    wire N__17893;
    wire N__17892;
    wire N__17891;
    wire N__17890;
    wire N__17887;
    wire N__17886;
    wire N__17885;
    wire N__17884;
    wire N__17881;
    wire N__17878;
    wire N__17875;
    wire N__17872;
    wire N__17869;
    wire N__17866;
    wire N__17859;
    wire N__17856;
    wire N__17855;
    wire N__17852;
    wire N__17841;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17827;
    wire N__17820;
    wire N__17817;
    wire N__17814;
    wire N__17811;
    wire N__17808;
    wire N__17801;
    wire N__17798;
    wire N__17793;
    wire N__17792;
    wire N__17791;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17773;
    wire N__17768;
    wire N__17763;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17748;
    wire N__17747;
    wire N__17744;
    wire N__17743;
    wire N__17736;
    wire N__17735;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17725;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17703;
    wire N__17702;
    wire N__17701;
    wire N__17700;
    wire N__17699;
    wire N__17698;
    wire N__17697;
    wire N__17696;
    wire N__17695;
    wire N__17694;
    wire N__17691;
    wire N__17686;
    wire N__17685;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17675;
    wire N__17666;
    wire N__17661;
    wire N__17652;
    wire N__17649;
    wire N__17646;
    wire N__17641;
    wire N__17634;
    wire N__17631;
    wire N__17628;
    wire N__17627;
    wire N__17626;
    wire N__17623;
    wire N__17618;
    wire N__17617;
    wire N__17616;
    wire N__17615;
    wire N__17610;
    wire N__17605;
    wire N__17602;
    wire N__17601;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17586;
    wire N__17577;
    wire N__17574;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17556;
    wire N__17555;
    wire N__17550;
    wire N__17549;
    wire N__17546;
    wire N__17545;
    wire N__17544;
    wire N__17541;
    wire N__17538;
    wire N__17533;
    wire N__17526;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17508;
    wire N__17507;
    wire N__17506;
    wire N__17505;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17493;
    wire N__17490;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17457;
    wire N__17456;
    wire N__17455;
    wire N__17454;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17439;
    wire N__17430;
    wire N__17427;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17409;
    wire N__17408;
    wire N__17403;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17395;
    wire N__17394;
    wire N__17393;
    wire N__17388;
    wire N__17381;
    wire N__17376;
    wire N__17375;
    wire N__17374;
    wire N__17371;
    wire N__17366;
    wire N__17363;
    wire N__17358;
    wire N__17357;
    wire N__17356;
    wire N__17355;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17341;
    wire N__17334;
    wire N__17331;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17292;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17280;
    wire N__17277;
    wire N__17276;
    wire N__17271;
    wire N__17268;
    wire N__17267;
    wire N__17264;
    wire N__17263;
    wire N__17262;
    wire N__17259;
    wire N__17252;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17237;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17217;
    wire N__17214;
    wire N__17213;
    wire N__17212;
    wire N__17207;
    wire N__17206;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17198;
    wire N__17197;
    wire N__17196;
    wire N__17195;
    wire N__17192;
    wire N__17191;
    wire N__17190;
    wire N__17187;
    wire N__17182;
    wire N__17175;
    wire N__17172;
    wire N__17167;
    wire N__17166;
    wire N__17165;
    wire N__17164;
    wire N__17163;
    wire N__17162;
    wire N__17161;
    wire N__17160;
    wire N__17159;
    wire N__17156;
    wire N__17155;
    wire N__17152;
    wire N__17147;
    wire N__17142;
    wire N__17133;
    wire N__17130;
    wire N__17129;
    wire N__17128;
    wire N__17125;
    wire N__17118;
    wire N__17115;
    wire N__17110;
    wire N__17107;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17091;
    wire N__17076;
    wire N__17075;
    wire N__17074;
    wire N__17071;
    wire N__17064;
    wire N__17061;
    wire N__17058;
    wire N__17055;
    wire N__17054;
    wire N__17053;
    wire N__17052;
    wire N__17051;
    wire N__17050;
    wire N__17049;
    wire N__17044;
    wire N__17043;
    wire N__17042;
    wire N__17041;
    wire N__17038;
    wire N__17037;
    wire N__17036;
    wire N__17027;
    wire N__17024;
    wire N__17023;
    wire N__17022;
    wire N__17019;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__16997;
    wire N__16992;
    wire N__16991;
    wire N__16990;
    wire N__16989;
    wire N__16988;
    wire N__16983;
    wire N__16980;
    wire N__16977;
    wire N__16972;
    wire N__16967;
    wire N__16956;
    wire N__16953;
    wire N__16952;
    wire N__16951;
    wire N__16948;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16932;
    wire N__16929;
    wire N__16928;
    wire N__16927;
    wire N__16926;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16908;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16890;
    wire N__16887;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16869;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16827;
    wire N__16826;
    wire N__16825;
    wire N__16824;
    wire N__16821;
    wire N__16820;
    wire N__16817;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16801;
    wire N__16800;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16785;
    wire N__16776;
    wire N__16773;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16755;
    wire N__16752;
    wire N__16749;
    wire N__16746;
    wire N__16743;
    wire N__16740;
    wire N__16737;
    wire N__16736;
    wire N__16731;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16719;
    wire N__16716;
    wire N__16713;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16677;
    wire N__16674;
    wire N__16671;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16647;
    wire N__16644;
    wire N__16643;
    wire N__16642;
    wire N__16641;
    wire N__16640;
    wire N__16639;
    wire N__16638;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16612;
    wire N__16609;
    wire N__16604;
    wire N__16599;
    wire N__16596;
    wire N__16589;
    wire N__16584;
    wire N__16581;
    wire N__16580;
    wire N__16577;
    wire N__16576;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16562;
    wire N__16561;
    wire N__16560;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16516;
    wire N__16507;
    wire N__16502;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16473;
    wire N__16470;
    wire N__16467;
    wire N__16466;
    wire N__16461;
    wire N__16458;
    wire N__16455;
    wire N__16452;
    wire N__16451;
    wire N__16448;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16358;
    wire N__16355;
    wire N__16354;
    wire N__16353;
    wire N__16352;
    wire N__16349;
    wire N__16340;
    wire N__16337;
    wire N__16332;
    wire N__16329;
    wire N__16328;
    wire N__16323;
    wire N__16320;
    wire N__16317;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16307;
    wire N__16306;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16293;
    wire N__16288;
    wire N__16281;
    wire N__16280;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16257;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16245;
    wire N__16242;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16230;
    wire N__16227;
    wire N__16224;
    wire N__16221;
    wire N__16218;
    wire N__16215;
    wire N__16212;
    wire N__16211;
    wire N__16210;
    wire N__16209;
    wire N__16208;
    wire N__16207;
    wire N__16206;
    wire N__16201;
    wire N__16198;
    wire N__16193;
    wire N__16192;
    wire N__16191;
    wire N__16186;
    wire N__16183;
    wire N__16178;
    wire N__16173;
    wire N__16164;
    wire N__16163;
    wire N__16162;
    wire N__16159;
    wire N__16158;
    wire N__16157;
    wire N__16156;
    wire N__16155;
    wire N__16154;
    wire N__16153;
    wire N__16152;
    wire N__16151;
    wire N__16150;
    wire N__16149;
    wire N__16148;
    wire N__16147;
    wire N__16146;
    wire N__16139;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16121;
    wire N__16118;
    wire N__16113;
    wire N__16108;
    wire N__16105;
    wire N__16104;
    wire N__16101;
    wire N__16100;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16088;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16067;
    wire N__16056;
    wire N__16051;
    wire N__16044;
    wire N__16041;
    wire N__16040;
    wire N__16035;
    wire N__16032;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16017;
    wire N__16014;
    wire N__16013;
    wire N__16012;
    wire N__16007;
    wire N__16004;
    wire N__15999;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15987;
    wire N__15984;
    wire N__15981;
    wire N__15978;
    wire N__15977;
    wire N__15976;
    wire N__15975;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15952;
    wire N__15949;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15924;
    wire N__15921;
    wire N__15920;
    wire N__15919;
    wire N__15916;
    wire N__15911;
    wire N__15908;
    wire N__15903;
    wire N__15902;
    wire N__15901;
    wire N__15900;
    wire N__15897;
    wire N__15896;
    wire N__15893;
    wire N__15892;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15880;
    wire N__15879;
    wire N__15878;
    wire N__15875;
    wire N__15870;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15853;
    wire N__15842;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15822;
    wire N__15819;
    wire N__15816;
    wire N__15813;
    wire N__15810;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15791;
    wire N__15790;
    wire N__15789;
    wire N__15788;
    wire N__15787;
    wire N__15784;
    wire N__15773;
    wire N__15770;
    wire N__15765;
    wire N__15764;
    wire N__15761;
    wire N__15756;
    wire N__15753;
    wire N__15750;
    wire N__15747;
    wire N__15744;
    wire N__15743;
    wire N__15742;
    wire N__15741;
    wire N__15738;
    wire N__15735;
    wire N__15730;
    wire N__15727;
    wire N__15720;
    wire N__15717;
    wire N__15714;
    wire N__15711;
    wire N__15708;
    wire N__15705;
    wire N__15702;
    wire N__15699;
    wire N__15698;
    wire N__15697;
    wire N__15696;
    wire N__15695;
    wire N__15692;
    wire N__15685;
    wire N__15682;
    wire N__15679;
    wire N__15672;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15657;
    wire N__15654;
    wire N__15651;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15641;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15624;
    wire N__15621;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15613;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15597;
    wire N__15596;
    wire N__15593;
    wire N__15590;
    wire N__15589;
    wire N__15588;
    wire N__15587;
    wire N__15576;
    wire N__15573;
    wire N__15570;
    wire N__15569;
    wire N__15568;
    wire N__15567;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15503;
    wire N__15500;
    wire N__15499;
    wire N__15498;
    wire N__15497;
    wire N__15496;
    wire N__15495;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15479;
    wire N__15474;
    wire N__15465;
    wire N__15462;
    wire N__15461;
    wire N__15460;
    wire N__15459;
    wire N__15458;
    wire N__15457;
    wire N__15456;
    wire N__15455;
    wire N__15452;
    wire N__15451;
    wire N__15450;
    wire N__15449;
    wire N__15448;
    wire N__15447;
    wire N__15444;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15430;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15411;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15399;
    wire N__15398;
    wire N__15395;
    wire N__15390;
    wire N__15387;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15367;
    wire N__15364;
    wire N__15361;
    wire N__15358;
    wire N__15355;
    wire N__15352;
    wire N__15347;
    wire N__15340;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15291;
    wire N__15288;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15246;
    wire N__15243;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15218;
    wire N__15215;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15198;
    wire N__15197;
    wire N__15196;
    wire N__15195;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15183;
    wire N__15182;
    wire N__15181;
    wire N__15180;
    wire N__15177;
    wire N__15172;
    wire N__15171;
    wire N__15170;
    wire N__15169;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15151;
    wire N__15142;
    wire N__15129;
    wire N__15128;
    wire N__15127;
    wire N__15126;
    wire N__15125;
    wire N__15124;
    wire N__15121;
    wire N__15120;
    wire N__15117;
    wire N__15116;
    wire N__15113;
    wire N__15108;
    wire N__15107;
    wire N__15106;
    wire N__15105;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15097;
    wire N__15096;
    wire N__15093;
    wire N__15092;
    wire N__15091;
    wire N__15088;
    wire N__15085;
    wire N__15084;
    wire N__15083;
    wire N__15080;
    wire N__15079;
    wire N__15076;
    wire N__15075;
    wire N__15074;
    wire N__15073;
    wire N__15072;
    wire N__15071;
    wire N__15070;
    wire N__15069;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15053;
    wire N__15042;
    wire N__15039;
    wire N__15036;
    wire N__15033;
    wire N__15030;
    wire N__15027;
    wire N__15024;
    wire N__15021;
    wire N__15018;
    wire N__15009;
    wire N__15004;
    wire N__14999;
    wire N__14994;
    wire N__14991;
    wire N__14964;
    wire N__14961;
    wire N__14958;
    wire N__14955;
    wire N__14952;
    wire N__14949;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14941;
    wire N__14940;
    wire N__14939;
    wire N__14938;
    wire N__14937;
    wire N__14936;
    wire N__14935;
    wire N__14932;
    wire N__14927;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14913;
    wire N__14910;
    wire N__14909;
    wire N__14904;
    wire N__14901;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14871;
    wire N__14860;
    wire N__14853;
    wire N__14852;
    wire N__14851;
    wire N__14850;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14836;
    wire N__14833;
    wire N__14830;
    wire N__14827;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14805;
    wire N__14802;
    wire N__14799;
    wire N__14796;
    wire N__14793;
    wire N__14790;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14778;
    wire N__14775;
    wire N__14772;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14745;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14727;
    wire N__14724;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14682;
    wire N__14679;
    wire N__14676;
    wire N__14673;
    wire N__14670;
    wire N__14667;
    wire N__14664;
    wire N__14661;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14653;
    wire N__14652;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14637;
    wire N__14636;
    wire N__14635;
    wire N__14634;
    wire N__14633;
    wire N__14632;
    wire N__14631;
    wire N__14630;
    wire N__14623;
    wire N__14612;
    wire N__14609;
    wire N__14604;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14592;
    wire N__14589;
    wire N__14584;
    wire N__14581;
    wire N__14574;
    wire N__14571;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14529;
    wire N__14528;
    wire N__14527;
    wire N__14526;
    wire N__14523;
    wire N__14522;
    wire N__14521;
    wire N__14520;
    wire N__14519;
    wire N__14518;
    wire N__14517;
    wire N__14516;
    wire N__14515;
    wire N__14514;
    wire N__14511;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14498;
    wire N__14493;
    wire N__14486;
    wire N__14483;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14475;
    wire N__14474;
    wire N__14471;
    wire N__14470;
    wire N__14469;
    wire N__14468;
    wire N__14465;
    wire N__14460;
    wire N__14455;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14433;
    wire N__14430;
    wire N__14425;
    wire N__14422;
    wire N__14419;
    wire N__14412;
    wire N__14407;
    wire N__14400;
    wire N__14385;
    wire N__14384;
    wire N__14383;
    wire N__14382;
    wire N__14381;
    wire N__14380;
    wire N__14375;
    wire N__14374;
    wire N__14373;
    wire N__14372;
    wire N__14371;
    wire N__14370;
    wire N__14367;
    wire N__14366;
    wire N__14361;
    wire N__14358;
    wire N__14355;
    wire N__14348;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14306;
    wire N__14299;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14274;
    wire N__14271;
    wire N__14268;
    wire N__14265;
    wire N__14262;
    wire N__14259;
    wire N__14256;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14238;
    wire N__14235;
    wire N__14232;
    wire N__14229;
    wire N__14226;
    wire N__14223;
    wire N__14220;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14208;
    wire N__14205;
    wire N__14202;
    wire N__14199;
    wire N__14196;
    wire N__14193;
    wire N__14190;
    wire N__14187;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14175;
    wire N__14172;
    wire N__14169;
    wire N__14166;
    wire N__14163;
    wire N__14160;
    wire N__14157;
    wire N__14154;
    wire N__14151;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14133;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14118;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14103;
    wire N__14100;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14088;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14073;
    wire N__14072;
    wire N__14069;
    wire N__14066;
    wire N__14063;
    wire N__14058;
    wire N__14055;
    wire N__14052;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14040;
    wire N__14037;
    wire N__14036;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14019;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14004;
    wire N__14001;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13968;
    wire N__13965;
    wire N__13962;
    wire N__13959;
    wire N__13956;
    wire N__13953;
    wire N__13950;
    wire N__13947;
    wire N__13944;
    wire N__13941;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13926;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13908;
    wire N__13905;
    wire N__13902;
    wire N__13899;
    wire N__13896;
    wire N__13893;
    wire N__13890;
    wire N__13889;
    wire N__13888;
    wire N__13887;
    wire N__13886;
    wire N__13877;
    wire N__13874;
    wire N__13869;
    wire N__13866;
    wire N__13865;
    wire N__13862;
    wire N__13861;
    wire N__13860;
    wire N__13859;
    wire N__13858;
    wire N__13857;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13843;
    wire N__13838;
    wire N__13827;
    wire N__13826;
    wire N__13823;
    wire N__13822;
    wire N__13821;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13803;
    wire N__13794;
    wire N__13793;
    wire N__13792;
    wire N__13791;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13781;
    wire N__13776;
    wire N__13767;
    wire N__13766;
    wire N__13765;
    wire N__13764;
    wire N__13757;
    wire N__13754;
    wire N__13749;
    wire N__13748;
    wire N__13747;
    wire N__13744;
    wire N__13739;
    wire N__13736;
    wire N__13731;
    wire N__13730;
    wire N__13727;
    wire N__13726;
    wire N__13725;
    wire N__13724;
    wire N__13723;
    wire N__13722;
    wire N__13721;
    wire N__13718;
    wire N__13717;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13703;
    wire N__13694;
    wire N__13691;
    wire N__13680;
    wire N__13677;
    wire N__13676;
    wire N__13675;
    wire N__13674;
    wire N__13673;
    wire N__13672;
    wire N__13671;
    wire N__13670;
    wire N__13669;
    wire N__13668;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13649;
    wire N__13646;
    wire N__13639;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13577;
    wire N__13572;
    wire N__13569;
    wire N__13566;
    wire N__13563;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13551;
    wire N__13550;
    wire N__13549;
    wire N__13548;
    wire N__13547;
    wire N__13546;
    wire N__13545;
    wire N__13542;
    wire N__13541;
    wire N__13538;
    wire N__13537;
    wire N__13534;
    wire N__13531;
    wire N__13524;
    wire N__13521;
    wire N__13518;
    wire N__13517;
    wire N__13510;
    wire N__13509;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13501;
    wire N__13498;
    wire N__13495;
    wire N__13494;
    wire N__13491;
    wire N__13488;
    wire N__13483;
    wire N__13478;
    wire N__13475;
    wire N__13470;
    wire N__13465;
    wire N__13462;
    wire N__13449;
    wire N__13448;
    wire N__13447;
    wire N__13446;
    wire N__13445;
    wire N__13444;
    wire N__13443;
    wire N__13442;
    wire N__13441;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13412;
    wire N__13411;
    wire N__13408;
    wire N__13405;
    wire N__13404;
    wire N__13401;
    wire N__13400;
    wire N__13399;
    wire N__13398;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13384;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13355;
    wire N__13354;
    wire N__13349;
    wire N__13346;
    wire N__13345;
    wire N__13342;
    wire N__13337;
    wire N__13332;
    wire N__13329;
    wire N__13326;
    wire N__13325;
    wire N__13324;
    wire N__13317;
    wire N__13314;
    wire N__13313;
    wire N__13310;
    wire N__13305;
    wire N__13302;
    wire N__13299;
    wire N__13296;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13269;
    wire N__13266;
    wire N__13263;
    wire N__13260;
    wire N__13259;
    wire N__13258;
    wire N__13255;
    wire N__13254;
    wire N__13251;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13224;
    wire N__13223;
    wire N__13220;
    wire N__13219;
    wire N__13216;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13172;
    wire N__13171;
    wire N__13170;
    wire N__13165;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13149;
    wire N__13148;
    wire N__13145;
    wire N__13144;
    wire N__13139;
    wire N__13136;
    wire N__13133;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13116;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13086;
    wire N__13083;
    wire N__13080;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13037;
    wire N__13034;
    wire N__13033;
    wire N__13032;
    wire N__13031;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13020;
    wire N__13019;
    wire N__13018;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13010;
    wire N__13007;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12993;
    wire N__12988;
    wire N__12985;
    wire N__12984;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12976;
    wire N__12975;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12946;
    wire N__12939;
    wire N__12924;
    wire N__12921;
    wire N__12918;
    wire N__12915;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12861;
    wire N__12860;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12830;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12816;
    wire N__12813;
    wire N__12810;
    wire N__12807;
    wire N__12806;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12791;
    wire N__12790;
    wire N__12789;
    wire N__12788;
    wire N__12787;
    wire N__12786;
    wire N__12785;
    wire N__12784;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12717;
    wire N__12714;
    wire N__12711;
    wire N__12708;
    wire N__12707;
    wire N__12702;
    wire N__12699;
    wire N__12698;
    wire N__12695;
    wire N__12692;
    wire N__12691;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12679;
    wire N__12672;
    wire N__12671;
    wire N__12668;
    wire N__12667;
    wire N__12666;
    wire N__12665;
    wire N__12660;
    wire N__12655;
    wire N__12652;
    wire N__12649;
    wire N__12646;
    wire N__12639;
    wire N__12638;
    wire N__12637;
    wire N__12636;
    wire N__12627;
    wire N__12626;
    wire N__12625;
    wire N__12622;
    wire N__12617;
    wire N__12616;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12570;
    wire N__12569;
    wire N__12568;
    wire N__12565;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12528;
    wire N__12525;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12513;
    wire N__12512;
    wire N__12511;
    wire N__12504;
    wire N__12501;
    wire N__12498;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12480;
    wire N__12479;
    wire N__12478;
    wire N__12477;
    wire N__12476;
    wire N__12473;
    wire N__12468;
    wire N__12463;
    wire N__12456;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12441;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12426;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12402;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12389;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12326;
    wire N__12325;
    wire N__12324;
    wire N__12323;
    wire N__12322;
    wire N__12321;
    wire N__12320;
    wire N__12317;
    wire N__12316;
    wire N__12315;
    wire N__12314;
    wire N__12313;
    wire N__12312;
    wire N__12311;
    wire N__12310;
    wire N__12299;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12281;
    wire N__12274;
    wire N__12269;
    wire N__12264;
    wire N__12255;
    wire N__12252;
    wire N__12249;
    wire N__12246;
    wire N__12243;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12219;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12198;
    wire N__12195;
    wire N__12192;
    wire N__12189;
    wire N__12188;
    wire N__12185;
    wire N__12182;
    wire N__12179;
    wire N__12176;
    wire N__12171;
    wire N__12168;
    wire N__12165;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12120;
    wire N__12117;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12089;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12081;
    wire N__12078;
    wire N__12073;
    wire N__12070;
    wire N__12067;
    wire N__12064;
    wire N__12061;
    wire N__12056;
    wire N__12053;
    wire N__12048;
    wire N__12047;
    wire N__12044;
    wire N__12043;
    wire N__12040;
    wire N__12037;
    wire N__12036;
    wire N__12035;
    wire N__12034;
    wire N__12031;
    wire N__12026;
    wire N__12023;
    wire N__12022;
    wire N__12021;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12007;
    wire N__12004;
    wire N__12001;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11975;
    wire N__11974;
    wire N__11973;
    wire N__11972;
    wire N__11971;
    wire N__11964;
    wire N__11963;
    wire N__11962;
    wire N__11959;
    wire N__11956;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11946;
    wire N__11943;
    wire N__11938;
    wire N__11935;
    wire N__11922;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11870;
    wire N__11869;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11847;
    wire N__11846;
    wire N__11845;
    wire N__11842;
    wire N__11841;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11830;
    wire N__11827;
    wire N__11824;
    wire N__11817;
    wire N__11814;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11792;
    wire N__11791;
    wire N__11788;
    wire N__11783;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11730;
    wire N__11727;
    wire N__11726;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11693;
    wire N__11692;
    wire N__11691;
    wire N__11690;
    wire N__11687;
    wire N__11678;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11664;
    wire N__11661;
    wire N__11660;
    wire N__11657;
    wire N__11656;
    wire N__11655;
    wire N__11652;
    wire N__11651;
    wire N__11648;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11628;
    wire N__11627;
    wire N__11624;
    wire N__11623;
    wire N__11622;
    wire N__11621;
    wire N__11618;
    wire N__11617;
    wire N__11612;
    wire N__11607;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11593;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11579;
    wire N__11576;
    wire N__11575;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire N__11553;
    wire N__11552;
    wire N__11549;
    wire N__11548;
    wire N__11547;
    wire N__11546;
    wire N__11545;
    wire N__11544;
    wire N__11541;
    wire N__11538;
    wire N__11529;
    wire N__11526;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11478;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11433;
    wire N__11432;
    wire N__11429;
    wire N__11426;
    wire N__11423;
    wire N__11420;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11337;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11307;
    wire N__11304;
    wire N__11303;
    wire N__11302;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11286;
    wire N__11283;
    wire N__11280;
    wire N__11277;
    wire N__11272;
    wire N__11269;
    wire N__11264;
    wire N__11261;
    wire N__11258;
    wire N__11253;
    wire N__11250;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11238;
    wire N__11235;
    wire N__11232;
    wire N__11231;
    wire N__11230;
    wire N__11225;
    wire N__11222;
    wire N__11217;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11193;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11169;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11151;
    wire N__11148;
    wire N__11145;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11124;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11108;
    wire N__11105;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11075;
    wire N__11074;
    wire N__11071;
    wire N__11066;
    wire N__11061;
    wire N__11060;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11025;
    wire N__11022;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10964;
    wire N__10959;
    wire N__10956;
    wire N__10953;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10941;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10923;
    wire N__10920;
    wire N__10917;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10902;
    wire N__10899;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10887;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10875;
    wire N__10872;
    wire N__10869;
    wire N__10866;
    wire N__10863;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10851;
    wire N__10848;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10832;
    wire N__10831;
    wire N__10830;
    wire N__10829;
    wire N__10828;
    wire N__10827;
    wire N__10824;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10804;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10788;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10761;
    wire N__10758;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10724;
    wire N__10723;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10715;
    wire N__10704;
    wire N__10701;
    wire N__10700;
    wire N__10697;
    wire N__10696;
    wire N__10695;
    wire N__10694;
    wire N__10693;
    wire N__10690;
    wire N__10685;
    wire N__10676;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10656;
    wire N__10653;
    wire N__10652;
    wire N__10651;
    wire N__10646;
    wire N__10643;
    wire N__10638;
    wire N__10635;
    wire N__10632;
    wire N__10631;
    wire N__10630;
    wire N__10629;
    wire N__10620;
    wire N__10617;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10589;
    wire N__10588;
    wire N__10585;
    wire N__10584;
    wire N__10581;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10556;
    wire N__10555;
    wire N__10554;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10538;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10512;
    wire N__10509;
    wire N__10506;
    wire N__10503;
    wire N__10500;
    wire N__10497;
    wire N__10494;
    wire N__10491;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10476;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10464;
    wire N__10463;
    wire N__10458;
    wire N__10455;
    wire N__10452;
    wire N__10451;
    wire N__10446;
    wire N__10445;
    wire N__10444;
    wire N__10441;
    wire N__10436;
    wire N__10431;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10419;
    wire N__10416;
    wire N__10413;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10405;
    wire N__10404;
    wire N__10403;
    wire N__10402;
    wire N__10401;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10389;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10356;
    wire N__10353;
    wire N__10350;
    wire N__10347;
    wire N__10344;
    wire N__10343;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10322;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10307;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10292;
    wire N__10289;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10269;
    wire N__10268;
    wire N__10267;
    wire N__10264;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10245;
    wire N__10242;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10206;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10182;
    wire N__10181;
    wire N__10180;
    wire N__10179;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10163;
    wire N__10162;
    wire N__10155;
    wire N__10152;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10140;
    wire N__10139;
    wire N__10136;
    wire N__10135;
    wire N__10134;
    wire N__10131;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10104;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10086;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10056;
    wire N__10053;
    wire N__10050;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10042;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10026;
    wire N__10023;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9965;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9946;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9930;
    wire N__9927;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9919;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9905;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9872;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9855;
    wire N__9854;
    wire N__9853;
    wire N__9852;
    wire N__9849;
    wire N__9840;
    wire N__9837;
    wire N__9834;
    wire N__9831;
    wire N__9830;
    wire N__9829;
    wire N__9828;
    wire N__9819;
    wire N__9816;
    wire N__9813;
    wire N__9810;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9800;
    wire N__9799;
    wire N__9796;
    wire N__9793;
    wire N__9792;
    wire N__9783;
    wire N__9780;
    wire N__9779;
    wire N__9778;
    wire N__9777;
    wire N__9768;
    wire N__9765;
    wire N__9762;
    wire N__9759;
    wire N__9756;
    wire N__9753;
    wire N__9752;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9735;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9725;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9708;
    wire N__9707;
    wire N__9706;
    wire N__9705;
    wire N__9702;
    wire N__9699;
    wire N__9694;
    wire N__9687;
    wire N__9684;
    wire N__9681;
    wire N__9680;
    wire N__9679;
    wire N__9678;
    wire N__9677;
    wire N__9674;
    wire N__9665;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9603;
    wire N__9602;
    wire N__9597;
    wire N__9594;
    wire N__9593;
    wire N__9590;
    wire N__9585;
    wire N__9582;
    wire N__9581;
    wire N__9578;
    wire N__9577;
    wire N__9574;
    wire N__9569;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9557;
    wire N__9556;
    wire N__9555;
    wire N__9554;
    wire N__9553;
    wire N__9552;
    wire N__9551;
    wire N__9544;
    wire N__9543;
    wire N__9532;
    wire N__9531;
    wire N__9530;
    wire N__9529;
    wire N__9528;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9506;
    wire N__9495;
    wire N__9492;
    wire N__9491;
    wire N__9490;
    wire N__9489;
    wire N__9488;
    wire N__9479;
    wire N__9478;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9466;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9446;
    wire N__9445;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9422;
    wire N__9419;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9390;
    wire N__9389;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9363;
    wire N__9360;
    wire N__9357;
    wire N__9354;
    wire N__9351;
    wire N__9348;
    wire N__9345;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9333;
    wire N__9330;
    wire N__9329;
    wire N__9328;
    wire N__9327;
    wire N__9322;
    wire N__9317;
    wire N__9312;
    wire N__9311;
    wire N__9308;
    wire N__9307;
    wire N__9306;
    wire N__9303;
    wire N__9298;
    wire N__9295;
    wire N__9288;
    wire N__9285;
    wire N__9284;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9261;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9251;
    wire N__9250;
    wire N__9249;
    wire N__9248;
    wire N__9247;
    wire N__9246;
    wire N__9245;
    wire N__9244;
    wire N__9243;
    wire N__9242;
    wire N__9241;
    wire N__9238;
    wire N__9231;
    wire N__9222;
    wire N__9213;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9197;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9171;
    wire N__9170;
    wire N__9169;
    wire N__9168;
    wire N__9167;
    wire N__9166;
    wire N__9165;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9157;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9143;
    wire N__9140;
    wire N__9131;
    wire N__9120;
    wire N__9119;
    wire N__9118;
    wire N__9117;
    wire N__9116;
    wire N__9113;
    wire N__9112;
    wire N__9111;
    wire N__9110;
    wire N__9107;
    wire N__9106;
    wire N__9105;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9082;
    wire N__9073;
    wire N__9066;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9056;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9039;
    wire N__9036;
    wire N__9033;
    wire N__9032;
    wire N__9029;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9016;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__9002;
    wire N__8999;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8979;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8965;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8939;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8922;
    wire N__8919;
    wire N__8916;
    wire N__8915;
    wire N__8912;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8823;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8783;
    wire N__8782;
    wire N__8781;
    wire N__8774;
    wire N__8771;
    wire N__8766;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8715;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8694;
    wire N__8691;
    wire N__8688;
    wire N__8687;
    wire N__8684;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8672;
    wire N__8671;
    wire N__8668;
    wire N__8667;
    wire N__8664;
    wire N__8657;
    wire N__8652;
    wire N__8651;
    wire N__8650;
    wire N__8649;
    wire N__8648;
    wire N__8645;
    wire N__8636;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8624;
    wire N__8619;
    wire N__8616;
    wire N__8615;
    wire N__8614;
    wire N__8607;
    wire N__8604;
    wire N__8603;
    wire N__8602;
    wire N__8599;
    wire N__8598;
    wire N__8597;
    wire N__8596;
    wire N__8591;
    wire N__8582;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8544;
    wire N__8541;
    wire N__8540;
    wire N__8537;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8523;
    wire N__8520;
    wire N__8517;
    wire N__8516;
    wire N__8511;
    wire N__8508;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8496;
    wire N__8495;
    wire N__8494;
    wire N__8491;
    wire N__8486;
    wire N__8481;
    wire N__8480;
    wire N__8477;
    wire N__8476;
    wire N__8473;
    wire N__8468;
    wire N__8463;
    wire N__8462;
    wire N__8459;
    wire N__8458;
    wire N__8457;
    wire N__8456;
    wire N__8455;
    wire N__8454;
    wire N__8451;
    wire N__8440;
    wire N__8435;
    wire N__8430;
    wire N__8429;
    wire N__8428;
    wire N__8421;
    wire N__8418;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8393;
    wire N__8388;
    wire N__8385;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8375;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8352;
    wire N__8349;
    wire N__8346;
    wire \latticehx1k_pll_inst.clk ;
    wire clk_in_c;
    wire GNDG0;
    wire VCCG0;
    wire bfn_1_1_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_ ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_0 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_0_cascade_ ;
    wire \buart.Z_tx.counter_RNIVE1P1_0_cascade_ ;
    wire \buart.Z_tx.un1_bitcount_c3_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire ufifo_utb_txdata_rdy_0_i_1_cascade_;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \buart.Z_tx.un1_bitcount_c2 ;
    wire ufifo_utb_txdata_rdy_0_i_1;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.counter_RNIVE1P1_0 ;
    wire ufifo_fifo_txdata_6;
    wire o_serial_data_c;
    wire \ufifo.fifo.fifo_txdata_7 ;
    wire N_366_cascade_;
    wire ufifo_utb_txdata_m0_7_cascade_;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire \ufifo.emitcrlf_fsm.cstate_ns_i_0_2_1_cascade_ ;
    wire \ufifo.N_323 ;
    wire \ufifo.emitcrlf_fsm.N_501_cascade_ ;
    wire \ufifo.emitcrlf_fsm.cstate_ns_i_0_0_1 ;
    wire bfn_1_6_0_;
    wire \ufifo.fifo.un1_wraddr_cry_0 ;
    wire \ufifo.fifo.un1_wraddr_cry_1 ;
    wire \ufifo.fifo.un1_wraddr_cry_2 ;
    wire \ufifo.fifo.un1_wraddr_cry_3 ;
    wire \ufifo.fifo.un1_wraddr_cry_4 ;
    wire \ufifo.fifo.un1_wraddr_cry_5 ;
    wire \ufifo.fifo.un1_wraddr_cry_6 ;
    wire \ufifo.fifo.un1_wraddr_cry_7 ;
    wire bfn_1_7_0_;
    wire ufifo_fifo_txdata_3;
    wire \buart.Z_tx.N_369_cascade_ ;
    wire ufifo_fifo_txdata_4;
    wire \buart.Z_tx.N_371_cascade_ ;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire N_366;
    wire ufifo_fifo_txdata_5;
    wire \buart.Z_tx.N_373_cascade_ ;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \buart.Z_tx.N_375 ;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire \buart.Z_tx.N_215_cascade_ ;
    wire N_257_cascade_;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0_cascade_ ;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire utb_txdata_1_cascade_;
    wire N_257;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire \buart.Z_tx.N_58 ;
    wire ufifo_emitcrlf_fsm_cstate_0;
    wire ufifo_emitcrlf_fsm_cstate_1;
    wire \ufifo.fifo.wraddrZ0Z_2 ;
    wire \ufifo.fifo.wraddrZ0Z_3 ;
    wire \ufifo.fifo.wraddrZ0Z_7 ;
    wire \ufifo.fifo.wraddrZ0Z_8 ;
    wire \ufifo.fifo.wraddrZ0Z_0 ;
    wire \ufifo.fifo.wraddrZ0Z_1 ;
    wire \ufifo.tx_fsm.N_358_cascade_ ;
    wire buart__tx_uart_busy_0;
    wire \ufifo.cstate_4 ;
    wire \ufifo.tx_fsm.N_394_cascade_ ;
    wire \ufifo.fifo.wraddrZ0Z_4 ;
    wire \ufifo.fifo.wraddrZ0Z_5 ;
    wire \ufifo.fifo.wraddrZ0Z_6 ;
    wire \ufifo.fifo.un1_emptyB_NE_0_cascade_ ;
    wire \ufifo.fifo.un1_emptyB_NE_3 ;
    wire \ufifo.fifo.un1_emptyB_NE_2 ;
    wire \ufifo.fifo.un1_emptyB_NE_4_cascade_ ;
    wire \ufifo.fifo.un1_emptyB_NE_1 ;
    wire \ufifo.emptyB_0_cascade_ ;
    wire \ufifo.tx_fsm.cstateZ0Z_5 ;
    wire \ufifo.tx_fsm.N_396_cascade_ ;
    wire \ufifo.tx_fsm.N_279 ;
    wire \ufifo.emptyB_0 ;
    wire \ufifo.tx_fsm.cstate_srsts_i_0_1_1_cascade_ ;
    wire \ufifo.tx_fsm.cstateZ0Z_1 ;
    wire \ufifo.fifo.fifo_txdata_2 ;
    wire \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0 ;
    wire \ufifo.sb_ram512x8_inst_RNILSN11_cascade_ ;
    wire utb_txdata_2;
    wire bfn_2_9_0_;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_rx.ser_clk ;
    wire \buart.Z_rx.N_76_i ;
    wire \Lab_UT.scdp.byteToEncrypt_7 ;
    wire \Lab_UT.scdp.prng_lfsr_7 ;
    wire \Lab_UT.scdp.prng_lfsr_15 ;
    wire \Lab_UT.scdp.lfsrInst.N_234_i_1_cascade_ ;
    wire uart_RXD;
    wire \Lab_UT.scdp.prng_lfsr_23 ;
    wire \resetGen.N_421_cascade_ ;
    wire \buart.Z_tx.N_554 ;
    wire \resetGen.N_267_cascade_ ;
    wire \resetGen.reset_countZ0Z_0 ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire \ufifo.popFifo ;
    wire \ufifo.fifo.rdaddrZ0Z_0 ;
    wire bfn_4_4_0_;
    wire \ufifo.fifo.rdaddrZ0Z_1 ;
    wire \ufifo.fifo.un1_rdaddr_cry_0 ;
    wire \ufifo.fifo.rdaddrZ0Z_2 ;
    wire \ufifo.fifo.un1_rdaddr_cry_1 ;
    wire \ufifo.fifo.rdaddrZ0Z_3 ;
    wire \ufifo.fifo.un1_rdaddr_cry_2 ;
    wire \ufifo.fifo.rdaddrZ0Z_4 ;
    wire \ufifo.fifo.un1_rdaddr_cry_3 ;
    wire \ufifo.fifo.rdaddrZ0Z_5 ;
    wire \ufifo.fifo.un1_rdaddr_cry_4 ;
    wire \ufifo.fifo.rdaddrZ0Z_6 ;
    wire \ufifo.fifo.un1_rdaddr_cry_5 ;
    wire \ufifo.fifo.rdaddrZ0Z_7 ;
    wire \ufifo.fifo.un1_rdaddr_cry_6 ;
    wire \ufifo.fifo.un1_rdaddr_cry_7 ;
    wire bfn_4_5_0_;
    wire \ufifo.fifo.rdaddrZ0Z_8 ;
    wire N_251;
    wire \ufifo.fifo.fifo_txdata_1 ;
    wire \ufifo.sb_ram512x8_inst_RNIKRN11 ;
    wire ufifo_fifo_txdata_rdy;
    wire \buart.Z_tx.N_278 ;
    wire \resetGen.N_274 ;
    wire \resetGen.N_421 ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire ufifo_tx_fsm_cstate_0;
    wire \ufifo.fifo.fifo_txdata_0 ;
    wire \Lab_UT.scdp.byteToEncrypt_0 ;
    wire \Lab_UT.scdp.byteToEncrypt_1 ;
    wire \Lab_UT.scdp.byteToEncrypt_2 ;
    wire \Lab_UT.scdp.b2a1.N_220_i_cascade_ ;
    wire \Lab_UT.scdp.b2a1.N_220_i ;
    wire \Lab_UT.scdp.N_282_cascade_ ;
    wire \Lab_UT.scdp.b2a1.N_293 ;
    wire \Lab_UT.scctrl.sccLdLFSR ;
    wire \Lab_UT.scctrl.EmsLoaded ;
    wire \Lab_UT.scctrl.EmsLoaded_cascade_ ;
    wire \Lab_UT.sccElsBitsLd_cascade_ ;
    wire \Lab_UT.scdp.lsBits_i_1_6 ;
    wire \Lab_UT.scdp.lsBitsD_6 ;
    wire \Lab_UT.scdp.N_282 ;
    wire \Lab_UT.scdp.byteToEncrypt_6 ;
    wire \Lab_UT.scdp.b2a0.N_238_i_cascade_ ;
    wire \Lab_UT.scdp.b2a0.N_238_i ;
    wire \Lab_UT.scdp.b2a0.N_227_i ;
    wire \Lab_UT.scdp.msBitsi.msBitsD_6 ;
    wire \Lab_UT.scdp.byteToEncrypt_5 ;
    wire \Lab_UT.scdp.b2a0.N_224_i ;
    wire \Lab_UT.scdp.msBitsi.msBitsD_0 ;
    wire \Lab_UT.scdp.lsBitsD_0 ;
    wire \Lab_UT.scdp.msBitsi.msBitsD_1 ;
    wire \Lab_UT.scdp.lsBitsD_1 ;
    wire \Lab_UT.scdp.msBitsi.N_43_cascade_ ;
    wire \ufifo.txdataDZ0Z_1 ;
    wire \Lab_UT.scdp.msBitsi.msBitsD_2 ;
    wire \Lab_UT.scdp.lsBitsD_2 ;
    wire \Lab_UT.scdp.msBitsi.msBitsD_4 ;
    wire \Lab_UT.scdp.lsBitsD_4 ;
    wire \Lab_UT.scdp.lsBitsi.lsBitsDZ0Z_5 ;
    wire \Lab_UT.scdp.N_332_i_1_cascade_ ;
    wire \ufifo.txdataDZ0Z_5 ;
    wire \Lab_UT.sccEmsBitsSl ;
    wire \Lab_UT.scdp.msBitsi.msBitsD_3 ;
    wire \Lab_UT.scdp.lsBitsD_3 ;
    wire \Lab_UT.scdp.g0_0_i_1_0 ;
    wire \Lab_UT.scdp.msBitsi.N_1915_0 ;
    wire \ufifo.txdataDZ0Z_3 ;
    wire \Lab_UT.scdp.msBitsi.N_1919_0 ;
    wire \ufifo.txdataDZ0Z_2 ;
    wire \Lab_UT.scdp.msBitsi.N_1917_0 ;
    wire \ufifo.txdataDZ0Z_4 ;
    wire \Lab_UT.scdp.N_552 ;
    wire \Lab_UT.scdp.N_228_i_0_cascade_ ;
    wire \Lab_UT.scdp.u0.byteToDecrypt_6 ;
    wire \Lab_UT.scdp.lfsrInst.N_234_i_0 ;
    wire \Lab_UT.scdp.g0_0_i_1 ;
    wire \Lab_UT.scdp.d2eData_3_0_1_cascade_ ;
    wire \Lab_UT.scdp.N_225_i_0 ;
    wire \Lab_UT.scdp.u1.g0_0_i_a5_0_2_cascade_ ;
    wire \Lab_UT.scdp.N_6 ;
    wire \Lab_UT.scdp.u1.g0_0_i_a5_0_2_0_cascade_ ;
    wire \Lab_UT.scdp.N_6_0 ;
    wire \Lab_UT.scdp.d2eData_3_0_a2_0_6 ;
    wire \Lab_UT.scdp.prng_lfsr_14 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30 ;
    wire \resetGen.N_243 ;
    wire \buart.bu_rx_data_i_2_4 ;
    wire \Lab_UT.scdp.msBitsi.q_esr_RNI679EZ0Z_6 ;
    wire \ufifo.txdataDZ0Z_6 ;
    wire \Lab_UT.scctrl.N_534 ;
    wire \Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0_cascade_ ;
    wire \Lab_UT.scctrl.N_415_0 ;
    wire \Lab_UT.scctrl.g1_0_0 ;
    wire \Lab_UT.scctrl.g1_0_2_cascade_ ;
    wire \Lab_UT.scctrl.next_state_0_0_2_cascade_ ;
    wire \ufifo.txDataValidDZ0 ;
    wire N_233_reti;
    wire \Lab_UT.scctrl.g1_0_1_0_cascade_ ;
    wire \Lab_UT.sccElsBitsLd ;
    wire \Lab_UT.scdp.sccElsBitsLd_0 ;
    wire \Lab_UT.scctrl.g1_0_1_cascade_ ;
    wire \Lab_UT.scdp.N_276 ;
    wire \Lab_UT.scdp.msBitsi.N_41 ;
    wire \ufifo.txdataDZ0Z_0 ;
    wire \Lab_UT.scctrl.N_46 ;
    wire \buart.Z_rx.sample_i_0_a2_0 ;
    wire \buart.Z_rx.N_230 ;
    wire \buart.Z_rx.N_230_cascade_ ;
    wire \Lab_UT.scdp.key0_7 ;
    wire \Lab_UT.scdp.key0_3 ;
    wire \Lab_UT.scdp.binVal_2_cascade_ ;
    wire \Lab_UT.scdp.N_73 ;
    wire \Lab_UT.scdp.N_73_cascade_ ;
    wire \Lab_UT.scctrl.delayload ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5 ;
    wire \Lab_UT.scdp.d2eData_3_5_cascade_ ;
    wire \Lab_UT.scdp.N_225_i_1 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21 ;
    wire \Lab_UT.scdp.u1.g0_0_i_a5_0_0_1_cascade_ ;
    wire \Lab_UT.scdp.u1.g0_0_i_a5_0_2_1 ;
    wire \Lab_UT.scdp.N_6_1 ;
    wire \Lab_UT.scdp.d2eData_3_0_3_cascade_ ;
    wire \Lab_UT.scdp.prng_lfsr_3 ;
    wire \Lab_UT.scdp.byteToEncrypt_3 ;
    wire \Lab_UT.scdp.d2eData_3_0_3 ;
    wire \Lab_UT.scdp.N_226_i ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19 ;
    wire \Lab_UT.scdp.d2eData_3_0_1 ;
    wire \Lab_UT.scdp.u1.byteToDecrypt_1 ;
    wire \Lab_UT.scdp.u1.N_539_cascade_ ;
    wire \Lab_UT.scdp.N_255_i ;
    wire \Lab_UT.scdp.N_228_i ;
    wire \Lab_UT.scdp.N_426_cascade_ ;
    wire \Lab_UT.scdp.q_RNI47LGA_1 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27 ;
    wire \Lab_UT.scdp.byteToEncrypt_4 ;
    wire \Lab_UT.scdp.b2a0.N_258_i ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1 ;
    wire \Lab_UT.scdp.d2eData_3_1_1 ;
    wire \Lab_UT.scdp.d2eData_3_0_a2_0_4 ;
    wire \Lab_UT.scdp.d2eData_3_0_a2_0_4_cascade_ ;
    wire \Lab_UT.scdp.N_246_i ;
    wire \Lab_UT.scdp.N_246_i_cascade_ ;
    wire \Lab_UT.scdp.u0.L4_tx_data_0_a2_1_6 ;
    wire \Lab_UT.scdp.N_256_i ;
    wire \Lab_UT.scdp.key0_2 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2 ;
    wire \Lab_UT.scdp.d2eData_3_2_cascade_ ;
    wire \Lab_UT.scdp.N_234_i ;
    wire \Lab_UT.scdp.byteToDecrypt_5 ;
    wire \Lab_UT.scdp.N_228_i_0 ;
    wire \Lab_UT.scdp.g0_0_i_0_cascade_ ;
    wire \Lab_UT.scdp.d2eData_3_5 ;
    wire \Lab_UT.scdp.g0_0_i_1_1 ;
    wire \Lab_UT.scctrl.g1_1_1_1_cascade_ ;
    wire \Lab_UT.scctrl.g2_0 ;
    wire \Lab_UT.scctrl.g1_3 ;
    wire \Lab_UT.scctrl.N_319_0 ;
    wire \Lab_UT.scctrl.N_414_0 ;
    wire \Lab_UT.scctrl.N_415_1_cascade_ ;
    wire \Lab_UT.scctrl.g1_0_0_0 ;
    wire \Lab_UT.scctrl.N_259i ;
    wire \Lab_UT.N_540i ;
    wire \Lab_UT.scctrl.N_266 ;
    wire \Lab_UT.scctrl.N_472_0 ;
    wire \Lab_UT.scctrl.N_241_reti ;
    wire \Lab_UT.scctrl.N_241_reti_cascade_ ;
    wire \Lab_UT.scctrl.N_263_0 ;
    wire \Lab_UT.scctrl.N_233_0 ;
    wire \Lab_UT.scctrl.N_351_1_0 ;
    wire \Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_5_1_cascade_ ;
    wire CONSTANT_ONE_NET_cascade_;
    wire \ufifo.sb_ram512x8_inst_RNIKTQ21 ;
    wire \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1Z0Z_0 ;
    wire N_368;
    wire utb_txdata_0;
    wire bfn_6_10_0_;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \buart.Z_rx.N_78 ;
    wire \Lab_UT.scctrl.N_418_0_cascade_ ;
    wire \Lab_UT.scctrl.g0_2 ;
    wire \Lab_UT.scctrl.g0_2_cascade_ ;
    wire \Lab_UT.scctrl.g1_1 ;
    wire \Lab_UT.scctrl.N_418_2_0_cascade_ ;
    wire \Lab_UT.scctrl.g1_1_2 ;
    wire \Lab_UT.scctrl.N_39_i_cascade_ ;
    wire \Lab_UT.scctrl.N_22_i_cascade_ ;
    wire \Lab_UT.state_1_ret_0_RNI9C1NH_0_cascade_ ;
    wire \Lab_UT.scdp.key3_5 ;
    wire \Lab_UT.state_1_ret_0_RNI9C1NH_0 ;
    wire \Lab_UT.scdp.key3_6 ;
    wire \Lab_UT.state_1_RNI6EDGH_0_2 ;
    wire \Lab_UT.scdp.key0_5 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0 ;
    wire \Lab_UT.scdp.d2eData_3_0_cascade_ ;
    wire \Lab_UT.scdp.N_262_i ;
    wire \Lab_UT.scdp.u1.g0_0_i_a5_0_0 ;
    wire \Lab_UT.scdp.d2eData_3_0 ;
    wire \Lab_UT.scdp.u1.byteToDecryptZ0Z_2 ;
    wire \Lab_UT.scdp.d2eData_3_2 ;
    wire \Lab_UT.scdp.u1.g0_0_i_a5_0_0_0 ;
    wire \Lab_UT.scdp.key0_6 ;
    wire \Lab_UT.scdp.prng_lfsr_6 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18 ;
    wire \Lab_UT.scdp.key0_4 ;
    wire \Lab_UT.scdp.prng_lfsr_4 ;
    wire \Lab_UT.scdp.key3_4 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28 ;
    wire \Lab_UT.scdp.prng_lfsr_11 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26 ;
    wire \Lab_UT.scdp.prng_lfsr_12 ;
    wire \Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9 ;
    wire \Lab_UT.sccLdLFSR_g ;
    wire \Lab_UT.scctrl.N_534_reti_cascade_ ;
    wire \Lab_UT.scctrl.N_266i ;
    wire bu_rx_data_2;
    wire \Lab_UT.N_540 ;
    wire \Lab_UT.scctrl.N_399_0 ;
    wire \Lab_UT.scctrl.sccEldByte_i_a2_0Z0Z_1 ;
    wire \Lab_UT.scctrl.g2 ;
    wire \Lab_UT.scctrl.g1_0_5 ;
    wire \Lab_UT.scctrl.next_state_1_0_2_cascade_ ;
    wire \Lab_UT.scctrl.N_444_0_cascade_ ;
    wire \Lab_UT.scctrl.N_319_1_0 ;
    wire \Lab_UT.scctrl.N_223_1_0_cascade_ ;
    wire \Lab_UT.scctrl.N_414_1_0 ;
    wire \Lab_UT.scctrl.N_444_0 ;
    wire \Lab_UT.scctrl.N_223_1_cascade_ ;
    wire \Lab_UT.scctrl.N_414_1_cascade_ ;
    wire \Lab_UT.scctrl.g1_0_2_0 ;
    wire \Lab_UT.scctrl.next_state_1_2_cascade_ ;
    wire \Lab_UT.scctrl.g0_0_i_0 ;
    wire \Lab_UT.scctrl.g0_0_i_1_cascade_ ;
    wire \Lab_UT.scctrl.g0_0_i_1_0_cascade_ ;
    wire \Lab_UT.scctrl.N_5_1 ;
    wire \Lab_UT.scctrl.g0_2_0_0_a3_1_1_cascade_ ;
    wire \Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0_cascade_ ;
    wire \Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0 ;
    wire \Lab_UT.scctrl.g0_i_o7_1_cascade_ ;
    wire \Lab_UT.scctrl.N_12_2_cascade_ ;
    wire bu_rx_data_i_2_3_rep1;
    wire \Lab_UT.scctrl.N_259 ;
    wire \Lab_UT.scctrl.g0_1_i_a8_0_1 ;
    wire \Lab_UT.scctrl.N_7_0 ;
    wire \Lab_UT.scctrl.N_10_0 ;
    wire \Lab_UT.scctrl.N_219 ;
    wire buart__rx_shifter_0_fast_1;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0_cascade_ ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0 ;
    wire buart__rx_shifter_2_fast_6;
    wire \Lab_UT.scctrl.N_444 ;
    wire bu_rx_data_i_2_fast_3;
    wire N_243_reti;
    wire \Lab_UT.scctrl.N_219i ;
    wire \Lab_UT.scctrl.N_271_0_0 ;
    wire \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_1_cascade_ ;
    wire buart__rx_shifter_0_fast_2;
    wire bu_rx_data_3;
    wire N_76_i_g;
    wire \buart.Z_rx.bitcountN11_15_i_0_o2_0_cascade_ ;
    wire \Lab_UT.scctrl.N_241 ;
    wire \Lab_UT.scctrl.g0_70_1_cascade_ ;
    wire \buart.Z_rx.N_80 ;
    wire \buart.Z_rx.bitcountZ0Z_0 ;
    wire \buart.Z_rx.bitcountZ0Z_3 ;
    wire \buart.Z_rx.bitcountZ0Z_2 ;
    wire buart__rx_N_86_i_0_o2_1_0;
    wire \Lab_UT.N_252 ;
    wire buart__rx_bitcount_4;
    wire buart__rx_N_86_i_0_o2_1_0_cascade_;
    wire buart__rx_bitcount_1;
    wire \Lab_UT.scctrl.r4.delay4 ;
    wire \Lab_UT.scctrl.delay3 ;
    wire \Lab_UT.scctrl.delay1 ;
    wire \Lab_UT.scctrl.delay2 ;
    wire \Lab_UT.scctrl.N_384 ;
    wire \Lab_UT.scctrl.N_385 ;
    wire \Lab_UT.scctrl.N_384_cascade_ ;
    wire \Lab_UT.N_100_i_cascade_ ;
    wire \Lab_UT.scdp.u2.N_100_i_0 ;
    wire \Lab_UT.scctrl.N_13_0_cascade_ ;
    wire \Lab_UT.scctrl.N_404_3_cascade_ ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_cascade_ ;
    wire \Lab_UT.scctrl.N_351 ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0 ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_0_0_cascade_ ;
    wire \Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_2 ;
    wire \Lab_UT.scctrl.N_6_2 ;
    wire \Lab_UT.scctrl.g0_8_1_0 ;
    wire \Lab_UT.scctrl.N_404_2 ;
    wire \Lab_UT.scctrl.g0_8_1_cascade_ ;
    wire \Lab_UT.scdp.key1_6 ;
    wire \Lab_UT.scdp.key1_7 ;
    wire \Lab_UT.scdp.key1_0 ;
    wire \Lab_UT.scdp.key1_3 ;
    wire \Lab_UT.scdp.key2_6 ;
    wire \Lab_UT.scdp.key2_4 ;
    wire \Lab_UT.scdp.key2_2 ;
    wire \Lab_UT.scdp.key1_2 ;
    wire \Lab_UT.scdp.key2_5 ;
    wire \Lab_UT.scdp.key1_4 ;
    wire \Lab_UT.scctrl.g1_0_4_cascade_ ;
    wire \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_3 ;
    wire \Lab_UT.scctrl.N_290_cascade_ ;
    wire \Lab_UT.scctrl.N_9_cascade_ ;
    wire \Lab_UT.scctrl.g0_9_0 ;
    wire \Lab_UT.scctrl.g0_1_2_0 ;
    wire \Lab_UT.scctrl.g3_cascade_ ;
    wire \Lab_UT.scctrl.g0_1_4 ;
    wire \Lab_UT.scctrl.next_state_rst_1_cascade_ ;
    wire \Lab_UT.scctrl.g0_i_0 ;
    wire \Lab_UT.scctrl.g3_0 ;
    wire \Lab_UT.scctrl.next_state_rst_0_7_cascade_ ;
    wire \Lab_UT.scctrl.N_10 ;
    wire \Lab_UT.scctrl.g0_1_i_0 ;
    wire \Lab_UT.scctrl.g0_1_i_2_cascade_ ;
    wire \Lab_UT.scctrl.g0_1_i_4 ;
    wire \Lab_UT.scctrl.next_state_rst_2_0 ;
    wire \Lab_UT.scctrl.G_24_i_a3_0_cascade_ ;
    wire \Lab_UT.scctrl.N_8 ;
    wire \Lab_UT.scctrl.N_290_2_cascade_ ;
    wire \Lab_UT.scctrl.N_8_3 ;
    wire \Lab_UT.scctrl.N_419_1 ;
    wire \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_2_3_cascade_ ;
    wire \Lab_UT.scctrl.g0_0_0 ;
    wire bu_rx_data_7;
    wire N_232;
    wire \Lab_UT.scctrl.g0_2_0 ;
    wire \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_1_3_cascade_ ;
    wire \Lab_UT.scctrl.next_state_0_0 ;
    wire \Lab_UT.scctrl.next_state_rst_cascade_ ;
    wire \Lab_UT.scctrl.state_i_1_0_rep2 ;
    wire \Lab_UT.scctrl.N_299_i_0_cascade_ ;
    wire \Lab_UT.scctrl.N_4 ;
    wire \Lab_UT.scctrl.N_240_reti ;
    wire \Lab_UT.scctrl.g0_2_0_0_a3_2_cascade_ ;
    wire \Lab_UT.scctrl.G_24_i_a3_3 ;
    wire \Lab_UT.scctrl.G_24_i_a3_5_cascade_ ;
    wire \Lab_UT.scctrl.G_24_i_a3_0_3 ;
    wire \Lab_UT.scctrl.G_24_i_a3_0_1 ;
    wire \Lab_UT.scctrl.N_15 ;
    wire \Lab_UT.scctrl.next_state_rst_0_3_tz_0 ;
    wire \Lab_UT.scctrl.g0_0_4_cascade_ ;
    wire \Lab_UT.scctrl.next_state_rst_4_1 ;
    wire \Lab_UT.scctrl.G_15_0_a10_1_2 ;
    wire \Lab_UT.scctrl.N_7 ;
    wire \Lab_UT.scctrl.g0_8_0_0 ;
    wire \Lab_UT.scctrl.N_223_0_0 ;
    wire \Lab_UT.scctrl.N_419_0_cascade_ ;
    wire \Lab_UT.scctrl.g1 ;
    wire \Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_0_3 ;
    wire \Lab_UT.scctrl.N_418_1 ;
    wire \Lab_UT.scctrl.g0_8_0_cascade_ ;
    wire \Lab_UT.scctrl.g0_8_2 ;
    wire \Lab_UT.scctrl.N_444_1 ;
    wire bu_rx_data_i_1_6;
    wire bu_rx_data_4;
    wire \Lab_UT.scctrl.G_24_i_a6_2_2_cascade_ ;
    wire \Lab_UT.scctrl.N_12_3 ;
    wire bu_rx_data_6;
    wire \Lab_UT.scctrl.N_241_i_0 ;
    wire \Lab_UT.scctrl.G_24_i_2_0 ;
    wire \Lab_UT.scctrl.G_24_i_a6_0_2 ;
    wire \Lab_UT.scctrl.N_5_2_cascade_ ;
    wire \Lab_UT.scctrl.next_state_rst_2_1 ;
    wire \Lab_UT.scctrl.G_24_i_1_0 ;
    wire \Lab_UT.scctrl.N_401_0 ;
    wire \Lab_UT.scctrl.N_9_0 ;
    wire \Lab_UT.scctrl.g0_i_2 ;
    wire \Lab_UT.scctrl.N_170_i_cascade_ ;
    wire \Lab_UT.scctrl.G_24_i_o6_0_0 ;
    wire \Lab_UT.scctrl.N_17_i_cascade_ ;
    wire \Lab_UT.scctrl.N_20_i_cascade_ ;
    wire \Lab_UT.scctrl.N_277 ;
    wire \Lab_UT.scctrl.N_277_cascade_ ;
    wire N_67;
    wire \Lab_UT.scctrl.N_355 ;
    wire \Lab_UT.scctrl.N_36 ;
    wire \Lab_UT.scctrl.N_27_i_cascade_ ;
    wire rst_i;
    wire \Lab_UT.scctrl.N_19 ;
    wire \Lab_UT.scctrl.N_415_2 ;
    wire \Lab_UT.scctrl.g1_2_0_cascade_ ;
    wire \Lab_UT.scctrl.next_stateZ0Z_2_cascade_ ;
    wire \Lab_UT.scctrl.next_state_rst_2 ;
    wire \Lab_UT.scctrl.next_stateZ0Z_2 ;
    wire \Lab_UT.scctrl.g1_1_1_0 ;
    wire \Lab_UT.scctrl.g1_2_0 ;
    wire \Lab_UT.scctrl.next_state_rst_4_3_cascade_ ;
    wire \Lab_UT.scctrl.N_290_0 ;
    wire \Lab_UT.scctrl.next_state_rst_4_5 ;
    wire \Lab_UT.scctrl.next_state_rst_4_4_cascade_ ;
    wire \Lab_UT.scctrl.N_290_1 ;
    wire \Lab_UT.scctrl.g0_1_0 ;
    wire \Lab_UT.scctrl.next_state_rst_1_3 ;
    wire \Lab_UT.scctrl.next_state_rst_4_2_cascade_ ;
    wire \Lab_UT.scctrl.N_290 ;
    wire \Lab_UT.scctrl.next_state_0_3 ;
    wire \Lab_UT.scctrl.N_418_2_cascade_ ;
    wire \Lab_UT.scctrl.g1_0 ;
    wire \Lab_UT.scctrl.N_418 ;
    wire \Lab_UT.scctrl.N_415 ;
    wire \Lab_UT.scctrl.state_ret_0_fastZ0 ;
    wire \Lab_UT.scctrl.state_ret_4_RNOZ0Z_10_cascade_ ;
    wire \Lab_UT.scctrl.state_ret_4_RNOZ0Z_6 ;
    wire \Lab_UT.scctrl.N_295 ;
    wire \Lab_UT.scctrl.N_295_cascade_ ;
    wire \Lab_UT.scctrl.N_40_i ;
    wire \Lab_UT.scctrl.N_487 ;
    wire \Lab_UT.scctrl.N_284 ;
    wire \Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0 ;
    wire \Lab_UT.scctrl.N_408_cascade_ ;
    wire \Lab_UT.scctrl.g0_i_a8_0_1_cascade_ ;
    wire \Lab_UT.scctrl.G_24_i_o7_0_0 ;
    wire \Lab_UT.scctrl.N_12_1_cascade_ ;
    wire \Lab_UT.scctrl.N_408 ;
    wire \Lab_UT.scctrl.next_state_rst_0_3_tz ;
    wire \Lab_UT.scctrl.next_state_rst_0_3_0_cascade_ ;
    wire rst_i_fast;
    wire \Lab_UT.scctrl.state_fast_3 ;
    wire \Lab_UT.scctrl.g0_0_0_0_cascade_ ;
    wire \Lab_UT.scctrl.g0_0_2_cascade_ ;
    wire \Lab_UT.scctrl.g0_0_3 ;
    wire buart__rx_shifter_1_fast_0;
    wire \Lab_UT.scctrl.N_408_0 ;
    wire \Lab_UT.scctrl.g2_0_0 ;
    wire \Lab_UT.scctrl.N_17 ;
    wire \Lab_UT.scctrl.N_240_i_0 ;
    wire bu_rx_data_i_1_5;
    wire \Lab_UT.scctrl.N_412_cascade_ ;
    wire \Lab_UT.scctrl.next_state_rst_0_1 ;
    wire \Lab_UT.scctrl.N_398i_i ;
    wire \Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0_0 ;
    wire \Lab_UT.scctrl.nibbleInZ0Z1 ;
    wire \Lab_UT.scctrl.N_69_cascade_ ;
    wire \Lab_UT.sccDnibble1En_cascade_ ;
    wire resetGen_rst_1_iso;
    wire \Lab_UT.scdp.u0.sccDnibble1En_0 ;
    wire \Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0dup_1 ;
    wire \Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93 ;
    wire \Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93_cascade_ ;
    wire \Lab_UT.scctrl.N_69_i ;
    wire \Lab_UT.scctrl.N_11 ;
    wire \Lab_UT.scctrl.next_state_rst ;
    wire \Lab_UT.scctrl.g0_9_a2_5_cascade_ ;
    wire \Lab_UT.scctrl.g1_1_0 ;
    wire \Lab_UT.scctrl.N_444_1_0 ;
    wire \Lab_UT.scctrl.g0_1_1 ;
    wire \Lab_UT.scctrl.g1_0_3_cascade_ ;
    wire \Lab_UT.scctrl.g1_2 ;
    wire \Lab_UT.scctrl.N_418_0_0 ;
    wire \Lab_UT.scctrl.g0_0 ;
    wire \Lab_UT.scctrl.g0_2_1 ;
    wire \Lab_UT.scctrl.g0_9_a2_2 ;
    wire \Lab_UT.scdp.byteToDecrypt_3 ;
    wire \Lab_UT.scdp.val_i_0_0_cascade_ ;
    wire \Lab_UT.scdp.a2b.N_280 ;
    wire bu_rx_data_0;
    wire \Lab_UT.scdp.N_378_cascade_ ;
    wire \Lab_UT.scdp.byteToDecrypt_4 ;
    wire \Lab_UT.scdp.val_i_0_0 ;
    wire \Lab_UT.scdp.N_378 ;
    wire \Lab_UT.scdp.u1.byteToDecryptZ0Z_0 ;
    wire \Lab_UT.scdp.a2b.val_0_tz_0_3 ;
    wire bu_rx_data_1;
    wire bu_rx_data_i_2_2;
    wire bu_rx_data_i_2_0;
    wire \Lab_UT.sccDnibble1En ;
    wire \Lab_UT.scdp.val_0_tz_3_cascade_ ;
    wire \Lab_UT.scdp.byteToDecrypt_7 ;
    wire \Lab_UT.scdp.key2_0 ;
    wire \Lab_UT.scdp.key2_1 ;
    wire \Lab_UT.scdp.key3_0 ;
    wire \Lab_UT.scdp.key3_1 ;
    wire \Lab_UT.scdp.binValD_2 ;
    wire \Lab_UT.scdp.key3_2 ;
    wire \Lab_UT.state_ret_12_RNIUVHQG_0 ;
    wire \Lab_UT.scdp.key3_3 ;
    wire \Lab_UT.scdp.val_0_tz_3 ;
    wire bu_rx_data_i_2_3;
    wire \buart.Z_rx.N_301 ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire buart__rx_hh_1;
    wire \buart.Z_rx.startbit ;
    wire \Lab_UT.scdp.binValD_0 ;
    wire \Lab_UT.scdp.key0_0 ;
    wire \Lab_UT.state_1_RNIO1RJH_0_2 ;
    wire \Lab_UT.scdp.key0_1 ;
    wire \Lab_UT.state_1_ret_3_RNI23U7H_0 ;
    wire \Lab_UT.scdp.key1_5 ;
    wire \Lab_UT.state_ret_RNIK5UKH_0 ;
    wire \Lab_UT.scdp.key2_3 ;
    wire \Lab_UT.scdp.binValD_1 ;
    wire \Lab_UT.state_ret_12_RNI2SEPG_0 ;
    wire \Lab_UT.scdp.key1_1 ;
    wire \Lab_UT.scdp.binVal_ValidD ;
    wire \Lab_UT.scdp.binValD_3 ;
    wire \Lab_UT.state_1_RNI2IGHH_0_0 ;
    wire \Lab_UT.scdp.key2_7 ;
    wire \Lab_UT.scctrl.state_i_1_0 ;
    wire \Lab_UT.scctrl.N_296_i_0 ;
    wire \Lab_UT.scctrl.next_state_RNO_1Z0Z_1 ;
    wire \Lab_UT.scctrl.N_319_cascade_ ;
    wire \Lab_UT.scctrl.next_state_rst_1_0 ;
    wire \Lab_UT.scctrl.N_414_cascade_ ;
    wire \Lab_UT.scctrl.next_state_rst_1_2 ;
    wire \Lab_UT.scctrl.N_319_1 ;
    wire \Lab_UT.scctrl.state_2_rep2 ;
    wire \Lab_UT.scctrl.N_7_1_cascade_ ;
    wire \Lab_UT.scctrl.G_18_i_a9_0_2 ;
    wire \Lab_UT.scctrl.G_18_i_1 ;
    wire \Lab_UT.scctrl.G_18_i_2_cascade_ ;
    wire \Lab_UT.scctrl.G_18_i_4_cascade_ ;
    wire \Lab_UT.scctrl.N_8_0_0 ;
    wire \Lab_UT.scctrl.g0_2_3_0 ;
    wire \Lab_UT.scctrl.g0_2_2_0 ;
    wire \Lab_UT.scctrl.next_state_2_0_cascade_ ;
    wire \Lab_UT.scctrl.N_260_i_0 ;
    wire \Lab_UT.scctrl.N_404_4 ;
    wire bu_rx_data_5;
    wire \Lab_UT.scctrl.g0_1_1_1 ;
    wire \Lab_UT.scctrl.g0_1_3 ;
    wire \Lab_UT.scctrl.next_state_rst_2_2 ;
    wire \Lab_UT.scctrl.N_13 ;
    wire \Lab_UT.scctrl.N_404_0 ;
    wire \Lab_UT.scctrl.N_5_3_cascade_ ;
    wire \Lab_UT.scctrl.N_12_0 ;
    wire \Lab_UT.scctrl.G_18_i_a9_0 ;
    wire \Lab_UT.scctrl.N_14_0 ;
    wire \Lab_UT.scctrl.stateZ0Z_2 ;
    wire \Lab_UT.scctrl.N_5 ;
    wire \Lab_UT.scctrl.N_21_0 ;
    wire \Lab_UT.scctrl.G_10_i_o7_0_cascade_ ;
    wire \Lab_UT.scctrl.G_24_i_a7_4_2 ;
    wire \Lab_UT.scctrl.G_24_i_1_cascade_ ;
    wire \Lab_UT.scctrl.N_13_2 ;
    wire \Lab_UT.scctrl.rst_retZ0 ;
    wire \Lab_UT.scctrl.state_i_2_2 ;
    wire \Lab_UT.scctrl.N_12_cascade_ ;
    wire \Lab_UT.scctrl.N_8_0 ;
    wire \Lab_UT.scctrl.g0_9_a2_4 ;
    wire \Lab_UT.scctrl.state_3_rep1 ;
    wire \Lab_UT.scctrl.g0_9_a3_0_0 ;
    wire \Lab_UT.scctrl.next_stateZ0Z_3 ;
    wire \Lab_UT.scctrl.next_state_0_1 ;
    wire \Lab_UT.scctrl.m90_i_o6_0_0_cascade_ ;
    wire \Lab_UT.scctrl.N_404_1 ;
    wire \Lab_UT.scctrl.N_401 ;
    wire \Lab_UT.scctrl.N_399 ;
    wire \Lab_UT.scctrl.g0_2_2_cascade_ ;
    wire \Lab_UT.scctrl.g0_2_3 ;
    wire \Lab_UT.scctrl.next_state_1_0_cascade_ ;
    wire \Lab_UT.scctrl.N_356_1_0 ;
    wire \Lab_UT.scctrl.g0_9_a2_1 ;
    wire \Lab_UT.scctrl.g0_2_3_1 ;
    wire \Lab_UT.scctrl.next_stateZ0Z_0 ;
    wire \Lab_UT.scctrl.g0_2_2_1 ;
    wire rst;
    wire \Lab_UT.scctrl.next_state_3_0 ;
    wire \Lab_UT.scctrl.next_stateZ0Z_1 ;
    wire \Lab_UT.scctrl.next_state_1_i_i_a2_1_0_1_cascade_ ;
    wire \Lab_UT.scctrl.next_state_rst_0_6 ;
    wire \Lab_UT.scctrl.N_398 ;
    wire \Lab_UT.scctrl.N_235_i_0 ;
    wire \Lab_UT.scctrl.N_240 ;
    wire \Lab_UT.scctrl.N_296 ;
    wire \Lab_UT.scctrl.state_1_ret_1_RNICEVZ0Z81 ;
    wire \Lab_UT.scctrl.N_72_i_cascade_ ;
    wire \Lab_UT.state_ret_11_RNI4RQC3_0 ;
    wire \Lab_UT.state_ret_11_RNI4RQC3_0_cascade_ ;
    wire N_74;
    wire \Lab_UT.sccDnibble2En ;
    wire \Lab_UT.scctrl.N_223 ;
    wire \Lab_UT.scctrl.stateZ0Z_0 ;
    wire \Lab_UT.scctrl.N_5_0 ;
    wire \Lab_UT.scctrl.G_10_i_a7_0_2 ;
    wire CONSTANT_ONE_NET;
    wire clk_g;
    wire \Lab_UT.scctrl.next_state_RNIN96CP1Z0Z_3 ;
    wire resetGen_rst_1_iso_g;
    wire \Lab_UT.scctrl.N_260 ;
    wire \Lab_UT.scctrl.N_235 ;
    wire N_55_i;
    wire \Lab_UT.scctrl.state_i_1_0_rep1 ;
    wire \Lab_UT.scctrl.state_2_rep1 ;
    wire \Lab_UT.scctrl.N_13_1 ;
    wire \Lab_UT.scctrl.G_10_i_1_cascade_ ;
    wire \Lab_UT.scctrl.state_fast_2 ;
    wire \Lab_UT.scctrl.state_i_1_fast_0 ;
    wire \Lab_UT.scctrl.next_state_0_2 ;
    wire rst_i_rep1;
    wire \Lab_UT.scctrl.N_21_cascade_ ;
    wire Lab_UT_scctrl_N_223_0;
    wire N_272;
    wire \Lab_UT.scctrl.G_15_0_1_cascade_ ;
    wire \Lab_UT.scctrl.stateZ0Z_3 ;
    wire \Lab_UT.scctrl.G_15_0_2 ;
    wire \Lab_UT.scctrl.state_i_2_3 ;
    wire N_21_1;
    wire \Lab_UT.scctrl.N_19_0 ;
    wire \Lab_UT.scctrl.N_8_1 ;
    wire \Lab_UT.scctrl.G_10_i_2 ;
    wire \Lab_UT.scctrl.G_24_i_0_cascade_ ;
    wire rst_ii;
    wire \Lab_UT.scctrl.G_24_i_2 ;
    wire \Lab_UT.scctrl.N_273 ;
    wire \Lab_UT.scctrl.N_261 ;
    wire \Lab_UT.scctrl.stateZ0Z_1 ;
    wire \Lab_UT.scctrl.N_8_2 ;
    wire \Lab_UT.N_245 ;
    wire N_245_i;
    wire _gnd_net_;

    defparam \ufifo.fifo.sb_ram512x8_inst_physical .WRITE_MODE=1;
    defparam \ufifo.fifo.sb_ram512x8_inst_physical .READ_MODE=1;
    SB_RAM40_4K \ufifo.fifo.sb_ram512x8_inst_physical  (
            .RDATA({dangling_wire_0,\ufifo.fifo.fifo_txdata_7 ,dangling_wire_1,ufifo_fifo_txdata_6,dangling_wire_2,ufifo_fifo_txdata_5,dangling_wire_3,ufifo_fifo_txdata_4,dangling_wire_4,ufifo_fifo_txdata_3,dangling_wire_5,\ufifo.fifo.fifo_txdata_2 ,dangling_wire_6,\ufifo.fifo.fifo_txdata_1 ,dangling_wire_7,\ufifo.fifo.fifo_txdata_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__10293,N__10326,N__9897,N__9927,N__9957,N__9990,N__10023,N__10056,N__10086}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__8979,N__9009,N__9399,N__9429,N__9456,N__9039,N__9066,N__8922,N__8949}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__11181,dangling_wire_31,N__10848,dangling_wire_32,N__10986,dangling_wire_33,N__10758,dangling_wire_34,N__11010,dangling_wire_35,N__10914,dangling_wire_36,N__11358}),
            .RCLKE(N__10140),
            .RCLK(N__21135),
            .RE(N__10130),
            .WCLKE(N__11302),
            .WCLK(N__21134),
            .WE(N__11307));
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\latticehx1k_pll_inst.clk ),
            .REFERENCECLK(N__8355),
            .RESETB(N__21192),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    IO_PAD led_obuf_4_iopad (
            .OE(N__23809),
            .DIN(N__23808),
            .DOUT(N__23807),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__23809),
            .PADOUT(N__23808),
            .PADIN(N__23807),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20541),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_1_iopad (
            .OE(N__23800),
            .DIN(N__23799),
            .DOUT(N__23798),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__23800),
            .PADOUT(N__23799),
            .PADIN(N__23798),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21588),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_3_iopad (
            .OE(N__23791),
            .DIN(N__23790),
            .DOUT(N__23789),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__23791),
            .PADOUT(N__23790),
            .PADIN(N__23789),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_0_iopad (
            .OE(N__23782),
            .DIN(N__23781),
            .DOUT(N__23780),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__23782),
            .PADOUT(N__23781),
            .PADIN(N__23780),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21633),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__23773),
            .DIN(N__23772),
            .DOUT(N__23771),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__23773),
            .PADOUT(N__23772),
            .PADIN(N__23771),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__21114),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__23764),
            .DIN(N__23763),
            .DOUT(N__23762),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__23764),
            .PADOUT(N__23763),
            .PADIN(N__23762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__23755),
            .DIN(N__23754),
            .DOUT(N__23753),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__23755),
            .PADOUT(N__23754),
            .PADIN(N__23753),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__23746),
            .DIN(N__23745),
            .DOUT(N__23744),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__23746),
            .PADOUT(N__23745),
            .PADIN(N__23744),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8562),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__23737),
            .DIN(N__23736),
            .DOUT(N__23735),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__23737),
            .PADOUT(N__23736),
            .PADIN(N__23735),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_2_iopad (
            .OE(N__23728),
            .DIN(N__23727),
            .DOUT(N__23726),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__23728),
            .PADOUT(N__23727),
            .PADIN(N__23726),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15525),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__5815 (
            .O(N__23709),
            .I(N__23701));
    CascadeMux I__5814 (
            .O(N__23708),
            .I(N__23698));
    CascadeMux I__5813 (
            .O(N__23707),
            .I(N__23692));
    InMux I__5812 (
            .O(N__23706),
            .I(N__23687));
    InMux I__5811 (
            .O(N__23705),
            .I(N__23676));
    InMux I__5810 (
            .O(N__23704),
            .I(N__23676));
    InMux I__5809 (
            .O(N__23701),
            .I(N__23676));
    InMux I__5808 (
            .O(N__23698),
            .I(N__23676));
    InMux I__5807 (
            .O(N__23697),
            .I(N__23676));
    InMux I__5806 (
            .O(N__23696),
            .I(N__23673));
    CascadeMux I__5805 (
            .O(N__23695),
            .I(N__23669));
    InMux I__5804 (
            .O(N__23692),
            .I(N__23663));
    InMux I__5803 (
            .O(N__23691),
            .I(N__23663));
    InMux I__5802 (
            .O(N__23690),
            .I(N__23660));
    LocalMux I__5801 (
            .O(N__23687),
            .I(N__23655));
    LocalMux I__5800 (
            .O(N__23676),
            .I(N__23655));
    LocalMux I__5799 (
            .O(N__23673),
            .I(N__23652));
    InMux I__5798 (
            .O(N__23672),
            .I(N__23649));
    InMux I__5797 (
            .O(N__23669),
            .I(N__23646));
    InMux I__5796 (
            .O(N__23668),
            .I(N__23643));
    LocalMux I__5795 (
            .O(N__23663),
            .I(N__23638));
    LocalMux I__5794 (
            .O(N__23660),
            .I(N__23638));
    Span4Mux_h I__5793 (
            .O(N__23655),
            .I(N__23635));
    Span4Mux_h I__5792 (
            .O(N__23652),
            .I(N__23630));
    LocalMux I__5791 (
            .O(N__23649),
            .I(N__23630));
    LocalMux I__5790 (
            .O(N__23646),
            .I(N__23625));
    LocalMux I__5789 (
            .O(N__23643),
            .I(N__23625));
    Span12Mux_s10_h I__5788 (
            .O(N__23638),
            .I(N__23622));
    Span4Mux_v I__5787 (
            .O(N__23635),
            .I(N__23619));
    Span4Mux_v I__5786 (
            .O(N__23630),
            .I(N__23614));
    Span4Mux_s1_h I__5785 (
            .O(N__23625),
            .I(N__23614));
    Odrv12 I__5784 (
            .O(N__23622),
            .I(\Lab_UT.scctrl.next_state_0_2 ));
    Odrv4 I__5783 (
            .O(N__23619),
            .I(\Lab_UT.scctrl.next_state_0_2 ));
    Odrv4 I__5782 (
            .O(N__23614),
            .I(\Lab_UT.scctrl.next_state_0_2 ));
    InMux I__5781 (
            .O(N__23607),
            .I(N__23601));
    InMux I__5780 (
            .O(N__23606),
            .I(N__23596));
    InMux I__5779 (
            .O(N__23605),
            .I(N__23593));
    InMux I__5778 (
            .O(N__23604),
            .I(N__23590));
    LocalMux I__5777 (
            .O(N__23601),
            .I(N__23586));
    InMux I__5776 (
            .O(N__23600),
            .I(N__23581));
    InMux I__5775 (
            .O(N__23599),
            .I(N__23581));
    LocalMux I__5774 (
            .O(N__23596),
            .I(N__23574));
    LocalMux I__5773 (
            .O(N__23593),
            .I(N__23574));
    LocalMux I__5772 (
            .O(N__23590),
            .I(N__23574));
    CascadeMux I__5771 (
            .O(N__23589),
            .I(N__23569));
    Span4Mux_v I__5770 (
            .O(N__23586),
            .I(N__23564));
    LocalMux I__5769 (
            .O(N__23581),
            .I(N__23564));
    Span4Mux_s3_h I__5768 (
            .O(N__23574),
            .I(N__23561));
    InMux I__5767 (
            .O(N__23573),
            .I(N__23558));
    InMux I__5766 (
            .O(N__23572),
            .I(N__23553));
    InMux I__5765 (
            .O(N__23569),
            .I(N__23553));
    Span4Mux_v I__5764 (
            .O(N__23564),
            .I(N__23550));
    Span4Mux_v I__5763 (
            .O(N__23561),
            .I(N__23547));
    LocalMux I__5762 (
            .O(N__23558),
            .I(N__23544));
    LocalMux I__5761 (
            .O(N__23553),
            .I(N__23535));
    Span4Mux_s3_h I__5760 (
            .O(N__23550),
            .I(N__23535));
    Span4Mux_s3_h I__5759 (
            .O(N__23547),
            .I(N__23535));
    Span4Mux_v I__5758 (
            .O(N__23544),
            .I(N__23535));
    Odrv4 I__5757 (
            .O(N__23535),
            .I(rst_i_rep1));
    CascadeMux I__5756 (
            .O(N__23532),
            .I(\Lab_UT.scctrl.N_21_cascade_ ));
    CascadeMux I__5755 (
            .O(N__23529),
            .I(N__23526));
    InMux I__5754 (
            .O(N__23526),
            .I(N__23520));
    InMux I__5753 (
            .O(N__23525),
            .I(N__23517));
    InMux I__5752 (
            .O(N__23524),
            .I(N__23514));
    CascadeMux I__5751 (
            .O(N__23523),
            .I(N__23510));
    LocalMux I__5750 (
            .O(N__23520),
            .I(N__23484));
    LocalMux I__5749 (
            .O(N__23517),
            .I(N__23481));
    LocalMux I__5748 (
            .O(N__23514),
            .I(N__23478));
    InMux I__5747 (
            .O(N__23513),
            .I(N__23475));
    InMux I__5746 (
            .O(N__23510),
            .I(N__23470));
    InMux I__5745 (
            .O(N__23509),
            .I(N__23470));
    InMux I__5744 (
            .O(N__23508),
            .I(N__23467));
    InMux I__5743 (
            .O(N__23507),
            .I(N__23464));
    InMux I__5742 (
            .O(N__23506),
            .I(N__23458));
    InMux I__5741 (
            .O(N__23505),
            .I(N__23458));
    InMux I__5740 (
            .O(N__23504),
            .I(N__23455));
    InMux I__5739 (
            .O(N__23503),
            .I(N__23449));
    CascadeMux I__5738 (
            .O(N__23502),
            .I(N__23445));
    CascadeMux I__5737 (
            .O(N__23501),
            .I(N__23435));
    CascadeMux I__5736 (
            .O(N__23500),
            .I(N__23430));
    CascadeMux I__5735 (
            .O(N__23499),
            .I(N__23427));
    CascadeMux I__5734 (
            .O(N__23498),
            .I(N__23422));
    InMux I__5733 (
            .O(N__23497),
            .I(N__23416));
    InMux I__5732 (
            .O(N__23496),
            .I(N__23416));
    InMux I__5731 (
            .O(N__23495),
            .I(N__23401));
    InMux I__5730 (
            .O(N__23494),
            .I(N__23401));
    InMux I__5729 (
            .O(N__23493),
            .I(N__23401));
    InMux I__5728 (
            .O(N__23492),
            .I(N__23401));
    InMux I__5727 (
            .O(N__23491),
            .I(N__23401));
    InMux I__5726 (
            .O(N__23490),
            .I(N__23401));
    InMux I__5725 (
            .O(N__23489),
            .I(N__23401));
    InMux I__5724 (
            .O(N__23488),
            .I(N__23398));
    CascadeMux I__5723 (
            .O(N__23487),
            .I(N__23395));
    Span4Mux_v I__5722 (
            .O(N__23484),
            .I(N__23381));
    Span4Mux_v I__5721 (
            .O(N__23481),
            .I(N__23381));
    Span4Mux_v I__5720 (
            .O(N__23478),
            .I(N__23381));
    LocalMux I__5719 (
            .O(N__23475),
            .I(N__23378));
    LocalMux I__5718 (
            .O(N__23470),
            .I(N__23373));
    LocalMux I__5717 (
            .O(N__23467),
            .I(N__23373));
    LocalMux I__5716 (
            .O(N__23464),
            .I(N__23370));
    InMux I__5715 (
            .O(N__23463),
            .I(N__23367));
    LocalMux I__5714 (
            .O(N__23458),
            .I(N__23362));
    LocalMux I__5713 (
            .O(N__23455),
            .I(N__23362));
    InMux I__5712 (
            .O(N__23454),
            .I(N__23359));
    InMux I__5711 (
            .O(N__23453),
            .I(N__23356));
    CascadeMux I__5710 (
            .O(N__23452),
            .I(N__23353));
    LocalMux I__5709 (
            .O(N__23449),
            .I(N__23345));
    InMux I__5708 (
            .O(N__23448),
            .I(N__23334));
    InMux I__5707 (
            .O(N__23445),
            .I(N__23334));
    InMux I__5706 (
            .O(N__23444),
            .I(N__23334));
    InMux I__5705 (
            .O(N__23443),
            .I(N__23334));
    InMux I__5704 (
            .O(N__23442),
            .I(N__23334));
    InMux I__5703 (
            .O(N__23441),
            .I(N__23323));
    InMux I__5702 (
            .O(N__23440),
            .I(N__23323));
    InMux I__5701 (
            .O(N__23439),
            .I(N__23323));
    InMux I__5700 (
            .O(N__23438),
            .I(N__23323));
    InMux I__5699 (
            .O(N__23435),
            .I(N__23323));
    InMux I__5698 (
            .O(N__23434),
            .I(N__23318));
    InMux I__5697 (
            .O(N__23433),
            .I(N__23318));
    InMux I__5696 (
            .O(N__23430),
            .I(N__23305));
    InMux I__5695 (
            .O(N__23427),
            .I(N__23305));
    InMux I__5694 (
            .O(N__23426),
            .I(N__23305));
    InMux I__5693 (
            .O(N__23425),
            .I(N__23305));
    InMux I__5692 (
            .O(N__23422),
            .I(N__23305));
    InMux I__5691 (
            .O(N__23421),
            .I(N__23305));
    LocalMux I__5690 (
            .O(N__23416),
            .I(N__23298));
    LocalMux I__5689 (
            .O(N__23401),
            .I(N__23298));
    LocalMux I__5688 (
            .O(N__23398),
            .I(N__23298));
    InMux I__5687 (
            .O(N__23395),
            .I(N__23293));
    InMux I__5686 (
            .O(N__23394),
            .I(N__23293));
    InMux I__5685 (
            .O(N__23393),
            .I(N__23280));
    InMux I__5684 (
            .O(N__23392),
            .I(N__23280));
    InMux I__5683 (
            .O(N__23391),
            .I(N__23280));
    InMux I__5682 (
            .O(N__23390),
            .I(N__23280));
    InMux I__5681 (
            .O(N__23389),
            .I(N__23280));
    InMux I__5680 (
            .O(N__23388),
            .I(N__23280));
    Span4Mux_v I__5679 (
            .O(N__23381),
            .I(N__23273));
    Span4Mux_v I__5678 (
            .O(N__23378),
            .I(N__23273));
    Span4Mux_v I__5677 (
            .O(N__23373),
            .I(N__23273));
    Span4Mux_h I__5676 (
            .O(N__23370),
            .I(N__23264));
    LocalMux I__5675 (
            .O(N__23367),
            .I(N__23264));
    Span4Mux_s3_h I__5674 (
            .O(N__23362),
            .I(N__23264));
    LocalMux I__5673 (
            .O(N__23359),
            .I(N__23264));
    LocalMux I__5672 (
            .O(N__23356),
            .I(N__23261));
    InMux I__5671 (
            .O(N__23353),
            .I(N__23252));
    InMux I__5670 (
            .O(N__23352),
            .I(N__23252));
    InMux I__5669 (
            .O(N__23351),
            .I(N__23252));
    InMux I__5668 (
            .O(N__23350),
            .I(N__23252));
    InMux I__5667 (
            .O(N__23349),
            .I(N__23247));
    InMux I__5666 (
            .O(N__23348),
            .I(N__23247));
    Span4Mux_v I__5665 (
            .O(N__23345),
            .I(N__23242));
    LocalMux I__5664 (
            .O(N__23334),
            .I(N__23242));
    LocalMux I__5663 (
            .O(N__23323),
            .I(N__23239));
    LocalMux I__5662 (
            .O(N__23318),
            .I(N__23230));
    LocalMux I__5661 (
            .O(N__23305),
            .I(N__23230));
    Span4Mux_v I__5660 (
            .O(N__23298),
            .I(N__23230));
    LocalMux I__5659 (
            .O(N__23293),
            .I(N__23230));
    LocalMux I__5658 (
            .O(N__23280),
            .I(Lab_UT_scctrl_N_223_0));
    Odrv4 I__5657 (
            .O(N__23273),
            .I(Lab_UT_scctrl_N_223_0));
    Odrv4 I__5656 (
            .O(N__23264),
            .I(Lab_UT_scctrl_N_223_0));
    Odrv12 I__5655 (
            .O(N__23261),
            .I(Lab_UT_scctrl_N_223_0));
    LocalMux I__5654 (
            .O(N__23252),
            .I(Lab_UT_scctrl_N_223_0));
    LocalMux I__5653 (
            .O(N__23247),
            .I(Lab_UT_scctrl_N_223_0));
    Odrv4 I__5652 (
            .O(N__23242),
            .I(Lab_UT_scctrl_N_223_0));
    Odrv12 I__5651 (
            .O(N__23239),
            .I(Lab_UT_scctrl_N_223_0));
    Odrv4 I__5650 (
            .O(N__23230),
            .I(Lab_UT_scctrl_N_223_0));
    InMux I__5649 (
            .O(N__23211),
            .I(N__23203));
    InMux I__5648 (
            .O(N__23210),
            .I(N__23203));
    InMux I__5647 (
            .O(N__23209),
            .I(N__23199));
    InMux I__5646 (
            .O(N__23208),
            .I(N__23192));
    LocalMux I__5645 (
            .O(N__23203),
            .I(N__23175));
    InMux I__5644 (
            .O(N__23202),
            .I(N__23172));
    LocalMux I__5643 (
            .O(N__23199),
            .I(N__23169));
    InMux I__5642 (
            .O(N__23198),
            .I(N__23166));
    InMux I__5641 (
            .O(N__23197),
            .I(N__23163));
    InMux I__5640 (
            .O(N__23196),
            .I(N__23157));
    InMux I__5639 (
            .O(N__23195),
            .I(N__23157));
    LocalMux I__5638 (
            .O(N__23192),
            .I(N__23154));
    InMux I__5637 (
            .O(N__23191),
            .I(N__23151));
    InMux I__5636 (
            .O(N__23190),
            .I(N__23144));
    InMux I__5635 (
            .O(N__23189),
            .I(N__23144));
    InMux I__5634 (
            .O(N__23188),
            .I(N__23141));
    InMux I__5633 (
            .O(N__23187),
            .I(N__23138));
    InMux I__5632 (
            .O(N__23186),
            .I(N__23129));
    InMux I__5631 (
            .O(N__23185),
            .I(N__23129));
    InMux I__5630 (
            .O(N__23184),
            .I(N__23129));
    InMux I__5629 (
            .O(N__23183),
            .I(N__23129));
    InMux I__5628 (
            .O(N__23182),
            .I(N__23123));
    InMux I__5627 (
            .O(N__23181),
            .I(N__23120));
    InMux I__5626 (
            .O(N__23180),
            .I(N__23112));
    InMux I__5625 (
            .O(N__23179),
            .I(N__23112));
    InMux I__5624 (
            .O(N__23178),
            .I(N__23109));
    Span4Mux_v I__5623 (
            .O(N__23175),
            .I(N__23105));
    LocalMux I__5622 (
            .O(N__23172),
            .I(N__23100));
    Span4Mux_v I__5621 (
            .O(N__23169),
            .I(N__23100));
    LocalMux I__5620 (
            .O(N__23166),
            .I(N__23097));
    LocalMux I__5619 (
            .O(N__23163),
            .I(N__23094));
    InMux I__5618 (
            .O(N__23162),
            .I(N__23091));
    LocalMux I__5617 (
            .O(N__23157),
            .I(N__23088));
    Span4Mux_s3_h I__5616 (
            .O(N__23154),
            .I(N__23083));
    LocalMux I__5615 (
            .O(N__23151),
            .I(N__23083));
    InMux I__5614 (
            .O(N__23150),
            .I(N__23080));
    InMux I__5613 (
            .O(N__23149),
            .I(N__23077));
    LocalMux I__5612 (
            .O(N__23144),
            .I(N__23074));
    LocalMux I__5611 (
            .O(N__23141),
            .I(N__23067));
    LocalMux I__5610 (
            .O(N__23138),
            .I(N__23067));
    LocalMux I__5609 (
            .O(N__23129),
            .I(N__23067));
    InMux I__5608 (
            .O(N__23128),
            .I(N__23064));
    InMux I__5607 (
            .O(N__23127),
            .I(N__23061));
    InMux I__5606 (
            .O(N__23126),
            .I(N__23058));
    LocalMux I__5605 (
            .O(N__23123),
            .I(N__23055));
    LocalMux I__5604 (
            .O(N__23120),
            .I(N__23052));
    InMux I__5603 (
            .O(N__23119),
            .I(N__23049));
    InMux I__5602 (
            .O(N__23118),
            .I(N__23044));
    InMux I__5601 (
            .O(N__23117),
            .I(N__23044));
    LocalMux I__5600 (
            .O(N__23112),
            .I(N__23039));
    LocalMux I__5599 (
            .O(N__23109),
            .I(N__23039));
    InMux I__5598 (
            .O(N__23108),
            .I(N__23036));
    Span4Mux_h I__5597 (
            .O(N__23105),
            .I(N__23023));
    Span4Mux_v I__5596 (
            .O(N__23100),
            .I(N__23023));
    Span4Mux_s2_h I__5595 (
            .O(N__23097),
            .I(N__23023));
    Span4Mux_v I__5594 (
            .O(N__23094),
            .I(N__23023));
    LocalMux I__5593 (
            .O(N__23091),
            .I(N__23023));
    Span4Mux_v I__5592 (
            .O(N__23088),
            .I(N__23023));
    Span4Mux_h I__5591 (
            .O(N__23083),
            .I(N__23010));
    LocalMux I__5590 (
            .O(N__23080),
            .I(N__23010));
    LocalMux I__5589 (
            .O(N__23077),
            .I(N__23010));
    Span4Mux_v I__5588 (
            .O(N__23074),
            .I(N__23010));
    Span4Mux_h I__5587 (
            .O(N__23067),
            .I(N__23010));
    LocalMux I__5586 (
            .O(N__23064),
            .I(N__23010));
    LocalMux I__5585 (
            .O(N__23061),
            .I(N__23005));
    LocalMux I__5584 (
            .O(N__23058),
            .I(N__23005));
    Span4Mux_v I__5583 (
            .O(N__23055),
            .I(N__23000));
    Span4Mux_s1_h I__5582 (
            .O(N__23052),
            .I(N__23000));
    LocalMux I__5581 (
            .O(N__23049),
            .I(N__22993));
    LocalMux I__5580 (
            .O(N__23044),
            .I(N__22993));
    Span4Mux_h I__5579 (
            .O(N__23039),
            .I(N__22993));
    LocalMux I__5578 (
            .O(N__23036),
            .I(N_272));
    Odrv4 I__5577 (
            .O(N__23023),
            .I(N_272));
    Odrv4 I__5576 (
            .O(N__23010),
            .I(N_272));
    Odrv4 I__5575 (
            .O(N__23005),
            .I(N_272));
    Odrv4 I__5574 (
            .O(N__23000),
            .I(N_272));
    Odrv4 I__5573 (
            .O(N__22993),
            .I(N_272));
    CascadeMux I__5572 (
            .O(N__22980),
            .I(\Lab_UT.scctrl.G_15_0_1_cascade_ ));
    CascadeMux I__5571 (
            .O(N__22977),
            .I(N__22972));
    InMux I__5570 (
            .O(N__22976),
            .I(N__22958));
    InMux I__5569 (
            .O(N__22975),
            .I(N__22954));
    InMux I__5568 (
            .O(N__22972),
            .I(N__22951));
    InMux I__5567 (
            .O(N__22971),
            .I(N__22948));
    InMux I__5566 (
            .O(N__22970),
            .I(N__22945));
    InMux I__5565 (
            .O(N__22969),
            .I(N__22941));
    InMux I__5564 (
            .O(N__22968),
            .I(N__22934));
    InMux I__5563 (
            .O(N__22967),
            .I(N__22934));
    InMux I__5562 (
            .O(N__22966),
            .I(N__22934));
    InMux I__5561 (
            .O(N__22965),
            .I(N__22927));
    InMux I__5560 (
            .O(N__22964),
            .I(N__22927));
    InMux I__5559 (
            .O(N__22963),
            .I(N__22927));
    InMux I__5558 (
            .O(N__22962),
            .I(N__22922));
    InMux I__5557 (
            .O(N__22961),
            .I(N__22922));
    LocalMux I__5556 (
            .O(N__22958),
            .I(N__22919));
    InMux I__5555 (
            .O(N__22957),
            .I(N__22915));
    LocalMux I__5554 (
            .O(N__22954),
            .I(N__22912));
    LocalMux I__5553 (
            .O(N__22951),
            .I(N__22909));
    LocalMux I__5552 (
            .O(N__22948),
            .I(N__22906));
    LocalMux I__5551 (
            .O(N__22945),
            .I(N__22903));
    InMux I__5550 (
            .O(N__22944),
            .I(N__22900));
    LocalMux I__5549 (
            .O(N__22941),
            .I(N__22895));
    LocalMux I__5548 (
            .O(N__22934),
            .I(N__22895));
    LocalMux I__5547 (
            .O(N__22927),
            .I(N__22892));
    LocalMux I__5546 (
            .O(N__22922),
            .I(N__22889));
    Sp12to4 I__5545 (
            .O(N__22919),
            .I(N__22885));
    InMux I__5544 (
            .O(N__22918),
            .I(N__22882));
    LocalMux I__5543 (
            .O(N__22915),
            .I(N__22877));
    Span4Mux_v I__5542 (
            .O(N__22912),
            .I(N__22877));
    Span4Mux_v I__5541 (
            .O(N__22909),
            .I(N__22872));
    Span4Mux_h I__5540 (
            .O(N__22906),
            .I(N__22872));
    Span4Mux_v I__5539 (
            .O(N__22903),
            .I(N__22865));
    LocalMux I__5538 (
            .O(N__22900),
            .I(N__22865));
    Span4Mux_v I__5537 (
            .O(N__22895),
            .I(N__22865));
    Span4Mux_s2_h I__5536 (
            .O(N__22892),
            .I(N__22860));
    Span4Mux_s2_h I__5535 (
            .O(N__22889),
            .I(N__22860));
    InMux I__5534 (
            .O(N__22888),
            .I(N__22857));
    Odrv12 I__5533 (
            .O(N__22885),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    LocalMux I__5532 (
            .O(N__22882),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    Odrv4 I__5531 (
            .O(N__22877),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    Odrv4 I__5530 (
            .O(N__22872),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    Odrv4 I__5529 (
            .O(N__22865),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    Odrv4 I__5528 (
            .O(N__22860),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    LocalMux I__5527 (
            .O(N__22857),
            .I(\Lab_UT.scctrl.stateZ0Z_3 ));
    InMux I__5526 (
            .O(N__22842),
            .I(N__22836));
    InMux I__5525 (
            .O(N__22841),
            .I(N__22836));
    LocalMux I__5524 (
            .O(N__22836),
            .I(N__22833));
    Odrv12 I__5523 (
            .O(N__22833),
            .I(\Lab_UT.scctrl.G_15_0_2 ));
    InMux I__5522 (
            .O(N__22830),
            .I(N__22816));
    InMux I__5521 (
            .O(N__22829),
            .I(N__22808));
    InMux I__5520 (
            .O(N__22828),
            .I(N__22808));
    InMux I__5519 (
            .O(N__22827),
            .I(N__22808));
    InMux I__5518 (
            .O(N__22826),
            .I(N__22805));
    InMux I__5517 (
            .O(N__22825),
            .I(N__22793));
    InMux I__5516 (
            .O(N__22824),
            .I(N__22793));
    InMux I__5515 (
            .O(N__22823),
            .I(N__22793));
    InMux I__5514 (
            .O(N__22822),
            .I(N__22793));
    InMux I__5513 (
            .O(N__22821),
            .I(N__22785));
    InMux I__5512 (
            .O(N__22820),
            .I(N__22782));
    InMux I__5511 (
            .O(N__22819),
            .I(N__22779));
    LocalMux I__5510 (
            .O(N__22816),
            .I(N__22776));
    InMux I__5509 (
            .O(N__22815),
            .I(N__22773));
    LocalMux I__5508 (
            .O(N__22808),
            .I(N__22770));
    LocalMux I__5507 (
            .O(N__22805),
            .I(N__22766));
    InMux I__5506 (
            .O(N__22804),
            .I(N__22761));
    InMux I__5505 (
            .O(N__22803),
            .I(N__22761));
    InMux I__5504 (
            .O(N__22802),
            .I(N__22758));
    LocalMux I__5503 (
            .O(N__22793),
            .I(N__22755));
    InMux I__5502 (
            .O(N__22792),
            .I(N__22752));
    InMux I__5501 (
            .O(N__22791),
            .I(N__22747));
    InMux I__5500 (
            .O(N__22790),
            .I(N__22747));
    InMux I__5499 (
            .O(N__22789),
            .I(N__22742));
    InMux I__5498 (
            .O(N__22788),
            .I(N__22742));
    LocalMux I__5497 (
            .O(N__22785),
            .I(N__22738));
    LocalMux I__5496 (
            .O(N__22782),
            .I(N__22733));
    LocalMux I__5495 (
            .O(N__22779),
            .I(N__22730));
    Span4Mux_s2_h I__5494 (
            .O(N__22776),
            .I(N__22723));
    LocalMux I__5493 (
            .O(N__22773),
            .I(N__22723));
    Span4Mux_h I__5492 (
            .O(N__22770),
            .I(N__22723));
    InMux I__5491 (
            .O(N__22769),
            .I(N__22720));
    Span4Mux_v I__5490 (
            .O(N__22766),
            .I(N__22717));
    LocalMux I__5489 (
            .O(N__22761),
            .I(N__22714));
    LocalMux I__5488 (
            .O(N__22758),
            .I(N__22707));
    Span4Mux_s3_v I__5487 (
            .O(N__22755),
            .I(N__22707));
    LocalMux I__5486 (
            .O(N__22752),
            .I(N__22707));
    LocalMux I__5485 (
            .O(N__22747),
            .I(N__22704));
    LocalMux I__5484 (
            .O(N__22742),
            .I(N__22701));
    InMux I__5483 (
            .O(N__22741),
            .I(N__22695));
    Span4Mux_s2_h I__5482 (
            .O(N__22738),
            .I(N__22692));
    InMux I__5481 (
            .O(N__22737),
            .I(N__22687));
    InMux I__5480 (
            .O(N__22736),
            .I(N__22687));
    Span12Mux_s6_h I__5479 (
            .O(N__22733),
            .I(N__22682));
    Span12Mux_s10_v I__5478 (
            .O(N__22730),
            .I(N__22682));
    Span4Mux_v I__5477 (
            .O(N__22723),
            .I(N__22679));
    LocalMux I__5476 (
            .O(N__22720),
            .I(N__22670));
    Span4Mux_s3_h I__5475 (
            .O(N__22717),
            .I(N__22670));
    Span4Mux_v I__5474 (
            .O(N__22714),
            .I(N__22670));
    Span4Mux_v I__5473 (
            .O(N__22707),
            .I(N__22670));
    Span4Mux_h I__5472 (
            .O(N__22704),
            .I(N__22665));
    Span4Mux_s2_h I__5471 (
            .O(N__22701),
            .I(N__22665));
    InMux I__5470 (
            .O(N__22700),
            .I(N__22658));
    InMux I__5469 (
            .O(N__22699),
            .I(N__22658));
    InMux I__5468 (
            .O(N__22698),
            .I(N__22658));
    LocalMux I__5467 (
            .O(N__22695),
            .I(\Lab_UT.scctrl.state_i_2_3 ));
    Odrv4 I__5466 (
            .O(N__22692),
            .I(\Lab_UT.scctrl.state_i_2_3 ));
    LocalMux I__5465 (
            .O(N__22687),
            .I(\Lab_UT.scctrl.state_i_2_3 ));
    Odrv12 I__5464 (
            .O(N__22682),
            .I(\Lab_UT.scctrl.state_i_2_3 ));
    Odrv4 I__5463 (
            .O(N__22679),
            .I(\Lab_UT.scctrl.state_i_2_3 ));
    Odrv4 I__5462 (
            .O(N__22670),
            .I(\Lab_UT.scctrl.state_i_2_3 ));
    Odrv4 I__5461 (
            .O(N__22665),
            .I(\Lab_UT.scctrl.state_i_2_3 ));
    LocalMux I__5460 (
            .O(N__22658),
            .I(\Lab_UT.scctrl.state_i_2_3 ));
    InMux I__5459 (
            .O(N__22641),
            .I(N__22638));
    LocalMux I__5458 (
            .O(N__22638),
            .I(N__22633));
    InMux I__5457 (
            .O(N__22637),
            .I(N__22630));
    InMux I__5456 (
            .O(N__22636),
            .I(N__22627));
    Span4Mux_h I__5455 (
            .O(N__22633),
            .I(N__22624));
    LocalMux I__5454 (
            .O(N__22630),
            .I(N_21_1));
    LocalMux I__5453 (
            .O(N__22627),
            .I(N_21_1));
    Odrv4 I__5452 (
            .O(N__22624),
            .I(N_21_1));
    CascadeMux I__5451 (
            .O(N__22617),
            .I(N__22614));
    InMux I__5450 (
            .O(N__22614),
            .I(N__22611));
    LocalMux I__5449 (
            .O(N__22611),
            .I(\Lab_UT.scctrl.N_19_0 ));
    InMux I__5448 (
            .O(N__22608),
            .I(N__22605));
    LocalMux I__5447 (
            .O(N__22605),
            .I(\Lab_UT.scctrl.N_8_1 ));
    InMux I__5446 (
            .O(N__22602),
            .I(N__22599));
    LocalMux I__5445 (
            .O(N__22599),
            .I(\Lab_UT.scctrl.G_10_i_2 ));
    CascadeMux I__5444 (
            .O(N__22596),
            .I(\Lab_UT.scctrl.G_24_i_0_cascade_ ));
    CascadeMux I__5443 (
            .O(N__22593),
            .I(N__22589));
    CascadeMux I__5442 (
            .O(N__22592),
            .I(N__22586));
    InMux I__5441 (
            .O(N__22589),
            .I(N__22577));
    InMux I__5440 (
            .O(N__22586),
            .I(N__22574));
    InMux I__5439 (
            .O(N__22585),
            .I(N__22571));
    InMux I__5438 (
            .O(N__22584),
            .I(N__22564));
    InMux I__5437 (
            .O(N__22583),
            .I(N__22564));
    InMux I__5436 (
            .O(N__22582),
            .I(N__22564));
    InMux I__5435 (
            .O(N__22581),
            .I(N__22558));
    InMux I__5434 (
            .O(N__22580),
            .I(N__22555));
    LocalMux I__5433 (
            .O(N__22577),
            .I(N__22552));
    LocalMux I__5432 (
            .O(N__22574),
            .I(N__22549));
    LocalMux I__5431 (
            .O(N__22571),
            .I(N__22543));
    LocalMux I__5430 (
            .O(N__22564),
            .I(N__22543));
    InMux I__5429 (
            .O(N__22563),
            .I(N__22531));
    InMux I__5428 (
            .O(N__22562),
            .I(N__22531));
    InMux I__5427 (
            .O(N__22561),
            .I(N__22531));
    LocalMux I__5426 (
            .O(N__22558),
            .I(N__22528));
    LocalMux I__5425 (
            .O(N__22555),
            .I(N__22525));
    Span4Mux_v I__5424 (
            .O(N__22552),
            .I(N__22520));
    Span4Mux_s3_h I__5423 (
            .O(N__22549),
            .I(N__22520));
    InMux I__5422 (
            .O(N__22548),
            .I(N__22517));
    Span4Mux_s3_h I__5421 (
            .O(N__22543),
            .I(N__22514));
    InMux I__5420 (
            .O(N__22542),
            .I(N__22511));
    InMux I__5419 (
            .O(N__22541),
            .I(N__22502));
    InMux I__5418 (
            .O(N__22540),
            .I(N__22502));
    InMux I__5417 (
            .O(N__22539),
            .I(N__22502));
    InMux I__5416 (
            .O(N__22538),
            .I(N__22502));
    LocalMux I__5415 (
            .O(N__22531),
            .I(N__22499));
    Span4Mux_h I__5414 (
            .O(N__22528),
            .I(N__22496));
    Span4Mux_v I__5413 (
            .O(N__22525),
            .I(N__22493));
    Span4Mux_h I__5412 (
            .O(N__22520),
            .I(N__22490));
    LocalMux I__5411 (
            .O(N__22517),
            .I(N__22485));
    Span4Mux_h I__5410 (
            .O(N__22514),
            .I(N__22485));
    LocalMux I__5409 (
            .O(N__22511),
            .I(rst_ii));
    LocalMux I__5408 (
            .O(N__22502),
            .I(rst_ii));
    Odrv12 I__5407 (
            .O(N__22499),
            .I(rst_ii));
    Odrv4 I__5406 (
            .O(N__22496),
            .I(rst_ii));
    Odrv4 I__5405 (
            .O(N__22493),
            .I(rst_ii));
    Odrv4 I__5404 (
            .O(N__22490),
            .I(rst_ii));
    Odrv4 I__5403 (
            .O(N__22485),
            .I(rst_ii));
    InMux I__5402 (
            .O(N__22470),
            .I(N__22467));
    LocalMux I__5401 (
            .O(N__22467),
            .I(\Lab_UT.scctrl.G_24_i_2 ));
    CascadeMux I__5400 (
            .O(N__22464),
            .I(N__22455));
    CascadeMux I__5399 (
            .O(N__22463),
            .I(N__22451));
    CascadeMux I__5398 (
            .O(N__22462),
            .I(N__22446));
    CascadeMux I__5397 (
            .O(N__22461),
            .I(N__22443));
    InMux I__5396 (
            .O(N__22460),
            .I(N__22437));
    InMux I__5395 (
            .O(N__22459),
            .I(N__22433));
    CascadeMux I__5394 (
            .O(N__22458),
            .I(N__22429));
    InMux I__5393 (
            .O(N__22455),
            .I(N__22425));
    CascadeMux I__5392 (
            .O(N__22454),
            .I(N__22421));
    InMux I__5391 (
            .O(N__22451),
            .I(N__22413));
    InMux I__5390 (
            .O(N__22450),
            .I(N__22413));
    InMux I__5389 (
            .O(N__22449),
            .I(N__22413));
    InMux I__5388 (
            .O(N__22446),
            .I(N__22410));
    InMux I__5387 (
            .O(N__22443),
            .I(N__22407));
    InMux I__5386 (
            .O(N__22442),
            .I(N__22404));
    CascadeMux I__5385 (
            .O(N__22441),
            .I(N__22401));
    CascadeMux I__5384 (
            .O(N__22440),
            .I(N__22397));
    LocalMux I__5383 (
            .O(N__22437),
            .I(N__22394));
    InMux I__5382 (
            .O(N__22436),
            .I(N__22391));
    LocalMux I__5381 (
            .O(N__22433),
            .I(N__22388));
    InMux I__5380 (
            .O(N__22432),
            .I(N__22383));
    InMux I__5379 (
            .O(N__22429),
            .I(N__22383));
    InMux I__5378 (
            .O(N__22428),
            .I(N__22380));
    LocalMux I__5377 (
            .O(N__22425),
            .I(N__22377));
    InMux I__5376 (
            .O(N__22424),
            .I(N__22372));
    InMux I__5375 (
            .O(N__22421),
            .I(N__22372));
    CascadeMux I__5374 (
            .O(N__22420),
            .I(N__22369));
    LocalMux I__5373 (
            .O(N__22413),
            .I(N__22366));
    LocalMux I__5372 (
            .O(N__22410),
            .I(N__22359));
    LocalMux I__5371 (
            .O(N__22407),
            .I(N__22359));
    LocalMux I__5370 (
            .O(N__22404),
            .I(N__22359));
    InMux I__5369 (
            .O(N__22401),
            .I(N__22356));
    InMux I__5368 (
            .O(N__22400),
            .I(N__22351));
    InMux I__5367 (
            .O(N__22397),
            .I(N__22351));
    Span4Mux_h I__5366 (
            .O(N__22394),
            .I(N__22342));
    LocalMux I__5365 (
            .O(N__22391),
            .I(N__22342));
    Span4Mux_s1_h I__5364 (
            .O(N__22388),
            .I(N__22342));
    LocalMux I__5363 (
            .O(N__22383),
            .I(N__22342));
    LocalMux I__5362 (
            .O(N__22380),
            .I(N__22339));
    Span4Mux_v I__5361 (
            .O(N__22377),
            .I(N__22334));
    LocalMux I__5360 (
            .O(N__22372),
            .I(N__22334));
    InMux I__5359 (
            .O(N__22369),
            .I(N__22331));
    Span4Mux_h I__5358 (
            .O(N__22366),
            .I(N__22326));
    Span4Mux_v I__5357 (
            .O(N__22359),
            .I(N__22326));
    LocalMux I__5356 (
            .O(N__22356),
            .I(N__22323));
    LocalMux I__5355 (
            .O(N__22351),
            .I(N__22316));
    Span4Mux_v I__5354 (
            .O(N__22342),
            .I(N__22316));
    Span4Mux_v I__5353 (
            .O(N__22339),
            .I(N__22316));
    Sp12to4 I__5352 (
            .O(N__22334),
            .I(N__22313));
    LocalMux I__5351 (
            .O(N__22331),
            .I(N__22308));
    Span4Mux_v I__5350 (
            .O(N__22326),
            .I(N__22308));
    Span4Mux_h I__5349 (
            .O(N__22323),
            .I(N__22303));
    Span4Mux_h I__5348 (
            .O(N__22316),
            .I(N__22303));
    Odrv12 I__5347 (
            .O(N__22313),
            .I(\Lab_UT.scctrl.N_273 ));
    Odrv4 I__5346 (
            .O(N__22308),
            .I(\Lab_UT.scctrl.N_273 ));
    Odrv4 I__5345 (
            .O(N__22303),
            .I(\Lab_UT.scctrl.N_273 ));
    InMux I__5344 (
            .O(N__22296),
            .I(N__22293));
    LocalMux I__5343 (
            .O(N__22293),
            .I(N__22281));
    InMux I__5342 (
            .O(N__22292),
            .I(N__22278));
    InMux I__5341 (
            .O(N__22291),
            .I(N__22275));
    InMux I__5340 (
            .O(N__22290),
            .I(N__22270));
    InMux I__5339 (
            .O(N__22289),
            .I(N__22270));
    InMux I__5338 (
            .O(N__22288),
            .I(N__22264));
    InMux I__5337 (
            .O(N__22287),
            .I(N__22261));
    InMux I__5336 (
            .O(N__22286),
            .I(N__22251));
    InMux I__5335 (
            .O(N__22285),
            .I(N__22251));
    InMux I__5334 (
            .O(N__22284),
            .I(N__22247));
    Span4Mux_v I__5333 (
            .O(N__22281),
            .I(N__22242));
    LocalMux I__5332 (
            .O(N__22278),
            .I(N__22242));
    LocalMux I__5331 (
            .O(N__22275),
            .I(N__22237));
    LocalMux I__5330 (
            .O(N__22270),
            .I(N__22237));
    InMux I__5329 (
            .O(N__22269),
            .I(N__22230));
    InMux I__5328 (
            .O(N__22268),
            .I(N__22230));
    InMux I__5327 (
            .O(N__22267),
            .I(N__22227));
    LocalMux I__5326 (
            .O(N__22264),
            .I(N__22224));
    LocalMux I__5325 (
            .O(N__22261),
            .I(N__22221));
    InMux I__5324 (
            .O(N__22260),
            .I(N__22210));
    InMux I__5323 (
            .O(N__22259),
            .I(N__22210));
    InMux I__5322 (
            .O(N__22258),
            .I(N__22210));
    InMux I__5321 (
            .O(N__22257),
            .I(N__22210));
    InMux I__5320 (
            .O(N__22256),
            .I(N__22210));
    LocalMux I__5319 (
            .O(N__22251),
            .I(N__22206));
    InMux I__5318 (
            .O(N__22250),
            .I(N__22203));
    LocalMux I__5317 (
            .O(N__22247),
            .I(N__22183));
    Span4Mux_h I__5316 (
            .O(N__22242),
            .I(N__22178));
    Span4Mux_s3_h I__5315 (
            .O(N__22237),
            .I(N__22178));
    InMux I__5314 (
            .O(N__22236),
            .I(N__22170));
    InMux I__5313 (
            .O(N__22235),
            .I(N__22170));
    LocalMux I__5312 (
            .O(N__22230),
            .I(N__22165));
    LocalMux I__5311 (
            .O(N__22227),
            .I(N__22165));
    Span4Mux_v I__5310 (
            .O(N__22224),
            .I(N__22158));
    Span4Mux_v I__5309 (
            .O(N__22221),
            .I(N__22158));
    LocalMux I__5308 (
            .O(N__22210),
            .I(N__22158));
    InMux I__5307 (
            .O(N__22209),
            .I(N__22155));
    Span4Mux_h I__5306 (
            .O(N__22206),
            .I(N__22150));
    LocalMux I__5305 (
            .O(N__22203),
            .I(N__22150));
    InMux I__5304 (
            .O(N__22202),
            .I(N__22141));
    InMux I__5303 (
            .O(N__22201),
            .I(N__22141));
    InMux I__5302 (
            .O(N__22200),
            .I(N__22141));
    InMux I__5301 (
            .O(N__22199),
            .I(N__22141));
    InMux I__5300 (
            .O(N__22198),
            .I(N__22134));
    InMux I__5299 (
            .O(N__22197),
            .I(N__22134));
    InMux I__5298 (
            .O(N__22196),
            .I(N__22134));
    InMux I__5297 (
            .O(N__22195),
            .I(N__22131));
    InMux I__5296 (
            .O(N__22194),
            .I(N__22126));
    InMux I__5295 (
            .O(N__22193),
            .I(N__22126));
    InMux I__5294 (
            .O(N__22192),
            .I(N__22123));
    InMux I__5293 (
            .O(N__22191),
            .I(N__22116));
    InMux I__5292 (
            .O(N__22190),
            .I(N__22116));
    InMux I__5291 (
            .O(N__22189),
            .I(N__22116));
    InMux I__5290 (
            .O(N__22188),
            .I(N__22109));
    InMux I__5289 (
            .O(N__22187),
            .I(N__22109));
    InMux I__5288 (
            .O(N__22186),
            .I(N__22109));
    Span4Mux_v I__5287 (
            .O(N__22183),
            .I(N__22104));
    Span4Mux_v I__5286 (
            .O(N__22178),
            .I(N__22104));
    InMux I__5285 (
            .O(N__22177),
            .I(N__22097));
    InMux I__5284 (
            .O(N__22176),
            .I(N__22097));
    InMux I__5283 (
            .O(N__22175),
            .I(N__22097));
    LocalMux I__5282 (
            .O(N__22170),
            .I(N__22090));
    Span4Mux_v I__5281 (
            .O(N__22165),
            .I(N__22090));
    Span4Mux_h I__5280 (
            .O(N__22158),
            .I(N__22090));
    LocalMux I__5279 (
            .O(N__22155),
            .I(N__22083));
    Span4Mux_v I__5278 (
            .O(N__22150),
            .I(N__22083));
    LocalMux I__5277 (
            .O(N__22141),
            .I(N__22083));
    LocalMux I__5276 (
            .O(N__22134),
            .I(N__22076));
    LocalMux I__5275 (
            .O(N__22131),
            .I(N__22076));
    LocalMux I__5274 (
            .O(N__22126),
            .I(N__22076));
    LocalMux I__5273 (
            .O(N__22123),
            .I(\Lab_UT.scctrl.N_261 ));
    LocalMux I__5272 (
            .O(N__22116),
            .I(\Lab_UT.scctrl.N_261 ));
    LocalMux I__5271 (
            .O(N__22109),
            .I(\Lab_UT.scctrl.N_261 ));
    Odrv4 I__5270 (
            .O(N__22104),
            .I(\Lab_UT.scctrl.N_261 ));
    LocalMux I__5269 (
            .O(N__22097),
            .I(\Lab_UT.scctrl.N_261 ));
    Odrv4 I__5268 (
            .O(N__22090),
            .I(\Lab_UT.scctrl.N_261 ));
    Odrv4 I__5267 (
            .O(N__22083),
            .I(\Lab_UT.scctrl.N_261 ));
    Odrv12 I__5266 (
            .O(N__22076),
            .I(\Lab_UT.scctrl.N_261 ));
    CascadeMux I__5265 (
            .O(N__22059),
            .I(N__22047));
    InMux I__5264 (
            .O(N__22058),
            .I(N__22038));
    InMux I__5263 (
            .O(N__22057),
            .I(N__22024));
    InMux I__5262 (
            .O(N__22056),
            .I(N__22019));
    InMux I__5261 (
            .O(N__22055),
            .I(N__22019));
    InMux I__5260 (
            .O(N__22054),
            .I(N__22016));
    InMux I__5259 (
            .O(N__22053),
            .I(N__22013));
    InMux I__5258 (
            .O(N__22052),
            .I(N__22010));
    InMux I__5257 (
            .O(N__22051),
            .I(N__22003));
    InMux I__5256 (
            .O(N__22050),
            .I(N__22003));
    InMux I__5255 (
            .O(N__22047),
            .I(N__22003));
    InMux I__5254 (
            .O(N__22046),
            .I(N__21998));
    InMux I__5253 (
            .O(N__22045),
            .I(N__21998));
    CascadeMux I__5252 (
            .O(N__22044),
            .I(N__21990));
    InMux I__5251 (
            .O(N__22043),
            .I(N__21986));
    InMux I__5250 (
            .O(N__22042),
            .I(N__21983));
    InMux I__5249 (
            .O(N__22041),
            .I(N__21980));
    LocalMux I__5248 (
            .O(N__22038),
            .I(N__21977));
    InMux I__5247 (
            .O(N__22037),
            .I(N__21966));
    InMux I__5246 (
            .O(N__22036),
            .I(N__21966));
    CascadeMux I__5245 (
            .O(N__22035),
            .I(N__21962));
    InMux I__5244 (
            .O(N__22034),
            .I(N__21957));
    InMux I__5243 (
            .O(N__22033),
            .I(N__21950));
    InMux I__5242 (
            .O(N__22032),
            .I(N__21950));
    InMux I__5241 (
            .O(N__22031),
            .I(N__21950));
    CascadeMux I__5240 (
            .O(N__22030),
            .I(N__21945));
    InMux I__5239 (
            .O(N__22029),
            .I(N__21938));
    InMux I__5238 (
            .O(N__22028),
            .I(N__21938));
    InMux I__5237 (
            .O(N__22027),
            .I(N__21938));
    LocalMux I__5236 (
            .O(N__22024),
            .I(N__21929));
    LocalMux I__5235 (
            .O(N__22019),
            .I(N__21929));
    LocalMux I__5234 (
            .O(N__22016),
            .I(N__21929));
    LocalMux I__5233 (
            .O(N__22013),
            .I(N__21929));
    LocalMux I__5232 (
            .O(N__22010),
            .I(N__21921));
    LocalMux I__5231 (
            .O(N__22003),
            .I(N__21921));
    LocalMux I__5230 (
            .O(N__21998),
            .I(N__21921));
    InMux I__5229 (
            .O(N__21997),
            .I(N__21910));
    InMux I__5228 (
            .O(N__21996),
            .I(N__21910));
    InMux I__5227 (
            .O(N__21995),
            .I(N__21910));
    InMux I__5226 (
            .O(N__21994),
            .I(N__21910));
    InMux I__5225 (
            .O(N__21993),
            .I(N__21910));
    InMux I__5224 (
            .O(N__21990),
            .I(N__21905));
    InMux I__5223 (
            .O(N__21989),
            .I(N__21905));
    LocalMux I__5222 (
            .O(N__21986),
            .I(N__21896));
    LocalMux I__5221 (
            .O(N__21983),
            .I(N__21896));
    LocalMux I__5220 (
            .O(N__21980),
            .I(N__21896));
    Span4Mux_s2_v I__5219 (
            .O(N__21977),
            .I(N__21896));
    InMux I__5218 (
            .O(N__21976),
            .I(N__21889));
    InMux I__5217 (
            .O(N__21975),
            .I(N__21889));
    InMux I__5216 (
            .O(N__21974),
            .I(N__21889));
    InMux I__5215 (
            .O(N__21973),
            .I(N__21882));
    InMux I__5214 (
            .O(N__21972),
            .I(N__21882));
    InMux I__5213 (
            .O(N__21971),
            .I(N__21882));
    LocalMux I__5212 (
            .O(N__21966),
            .I(N__21879));
    InMux I__5211 (
            .O(N__21965),
            .I(N__21876));
    InMux I__5210 (
            .O(N__21962),
            .I(N__21867));
    InMux I__5209 (
            .O(N__21961),
            .I(N__21867));
    InMux I__5208 (
            .O(N__21960),
            .I(N__21864));
    LocalMux I__5207 (
            .O(N__21957),
            .I(N__21859));
    LocalMux I__5206 (
            .O(N__21950),
            .I(N__21859));
    CascadeMux I__5205 (
            .O(N__21949),
            .I(N__21855));
    InMux I__5204 (
            .O(N__21948),
            .I(N__21850));
    InMux I__5203 (
            .O(N__21945),
            .I(N__21847));
    LocalMux I__5202 (
            .O(N__21938),
            .I(N__21842));
    Span4Mux_v I__5201 (
            .O(N__21929),
            .I(N__21842));
    InMux I__5200 (
            .O(N__21928),
            .I(N__21839));
    Span4Mux_v I__5199 (
            .O(N__21921),
            .I(N__21836));
    LocalMux I__5198 (
            .O(N__21910),
            .I(N__21831));
    LocalMux I__5197 (
            .O(N__21905),
            .I(N__21831));
    Span4Mux_v I__5196 (
            .O(N__21896),
            .I(N__21828));
    LocalMux I__5195 (
            .O(N__21889),
            .I(N__21819));
    LocalMux I__5194 (
            .O(N__21882),
            .I(N__21819));
    Span4Mux_h I__5193 (
            .O(N__21879),
            .I(N__21819));
    LocalMux I__5192 (
            .O(N__21876),
            .I(N__21819));
    InMux I__5191 (
            .O(N__21875),
            .I(N__21809));
    InMux I__5190 (
            .O(N__21874),
            .I(N__21809));
    InMux I__5189 (
            .O(N__21873),
            .I(N__21809));
    InMux I__5188 (
            .O(N__21872),
            .I(N__21806));
    LocalMux I__5187 (
            .O(N__21867),
            .I(N__21803));
    LocalMux I__5186 (
            .O(N__21864),
            .I(N__21798));
    Span4Mux_v I__5185 (
            .O(N__21859),
            .I(N__21798));
    InMux I__5184 (
            .O(N__21858),
            .I(N__21795));
    InMux I__5183 (
            .O(N__21855),
            .I(N__21792));
    InMux I__5182 (
            .O(N__21854),
            .I(N__21787));
    InMux I__5181 (
            .O(N__21853),
            .I(N__21787));
    LocalMux I__5180 (
            .O(N__21850),
            .I(N__21780));
    LocalMux I__5179 (
            .O(N__21847),
            .I(N__21780));
    Span4Mux_h I__5178 (
            .O(N__21842),
            .I(N__21780));
    LocalMux I__5177 (
            .O(N__21839),
            .I(N__21775));
    Span4Mux_h I__5176 (
            .O(N__21836),
            .I(N__21775));
    Span4Mux_v I__5175 (
            .O(N__21831),
            .I(N__21768));
    Span4Mux_h I__5174 (
            .O(N__21828),
            .I(N__21768));
    Span4Mux_v I__5173 (
            .O(N__21819),
            .I(N__21768));
    InMux I__5172 (
            .O(N__21818),
            .I(N__21761));
    InMux I__5171 (
            .O(N__21817),
            .I(N__21761));
    InMux I__5170 (
            .O(N__21816),
            .I(N__21761));
    LocalMux I__5169 (
            .O(N__21809),
            .I(N__21758));
    LocalMux I__5168 (
            .O(N__21806),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    Odrv4 I__5167 (
            .O(N__21803),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    Odrv4 I__5166 (
            .O(N__21798),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    LocalMux I__5165 (
            .O(N__21795),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    LocalMux I__5164 (
            .O(N__21792),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    LocalMux I__5163 (
            .O(N__21787),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    Odrv4 I__5162 (
            .O(N__21780),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    Odrv4 I__5161 (
            .O(N__21775),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    Odrv4 I__5160 (
            .O(N__21768),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    LocalMux I__5159 (
            .O(N__21761),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    Odrv12 I__5158 (
            .O(N__21758),
            .I(\Lab_UT.scctrl.stateZ0Z_1 ));
    InMux I__5157 (
            .O(N__21735),
            .I(N__21732));
    LocalMux I__5156 (
            .O(N__21732),
            .I(\Lab_UT.scctrl.N_8_2 ));
    CascadeMux I__5155 (
            .O(N__21729),
            .I(N__21725));
    CascadeMux I__5154 (
            .O(N__21728),
            .I(N__21718));
    InMux I__5153 (
            .O(N__21725),
            .I(N__21714));
    InMux I__5152 (
            .O(N__21724),
            .I(N__21711));
    CascadeMux I__5151 (
            .O(N__21723),
            .I(N__21703));
    InMux I__5150 (
            .O(N__21722),
            .I(N__21700));
    InMux I__5149 (
            .O(N__21721),
            .I(N__21697));
    InMux I__5148 (
            .O(N__21718),
            .I(N__21692));
    InMux I__5147 (
            .O(N__21717),
            .I(N__21692));
    LocalMux I__5146 (
            .O(N__21714),
            .I(N__21687));
    LocalMux I__5145 (
            .O(N__21711),
            .I(N__21687));
    InMux I__5144 (
            .O(N__21710),
            .I(N__21682));
    InMux I__5143 (
            .O(N__21709),
            .I(N__21682));
    InMux I__5142 (
            .O(N__21708),
            .I(N__21677));
    InMux I__5141 (
            .O(N__21707),
            .I(N__21677));
    InMux I__5140 (
            .O(N__21706),
            .I(N__21672));
    InMux I__5139 (
            .O(N__21703),
            .I(N__21672));
    LocalMux I__5138 (
            .O(N__21700),
            .I(N__21669));
    LocalMux I__5137 (
            .O(N__21697),
            .I(N__21666));
    LocalMux I__5136 (
            .O(N__21692),
            .I(N__21663));
    Span4Mux_v I__5135 (
            .O(N__21687),
            .I(N__21660));
    LocalMux I__5134 (
            .O(N__21682),
            .I(N__21653));
    LocalMux I__5133 (
            .O(N__21677),
            .I(N__21653));
    LocalMux I__5132 (
            .O(N__21672),
            .I(N__21653));
    Span4Mux_v I__5131 (
            .O(N__21669),
            .I(N__21650));
    Span4Mux_h I__5130 (
            .O(N__21666),
            .I(N__21645));
    Span4Mux_v I__5129 (
            .O(N__21663),
            .I(N__21645));
    Sp12to4 I__5128 (
            .O(N__21660),
            .I(N__21640));
    Span12Mux_s8_v I__5127 (
            .O(N__21653),
            .I(N__21640));
    Odrv4 I__5126 (
            .O(N__21650),
            .I(\Lab_UT.N_245 ));
    Odrv4 I__5125 (
            .O(N__21645),
            .I(\Lab_UT.N_245 ));
    Odrv12 I__5124 (
            .O(N__21640),
            .I(\Lab_UT.N_245 ));
    IoInMux I__5123 (
            .O(N__21633),
            .I(N__21630));
    LocalMux I__5122 (
            .O(N__21630),
            .I(N_245_i));
    CascadeMux I__5121 (
            .O(N__21627),
            .I(\Lab_UT.scctrl.N_72_i_cascade_ ));
    InMux I__5120 (
            .O(N__21624),
            .I(N__21615));
    InMux I__5119 (
            .O(N__21623),
            .I(N__21615));
    InMux I__5118 (
            .O(N__21622),
            .I(N__21615));
    LocalMux I__5117 (
            .O(N__21615),
            .I(N__21612));
    Span4Mux_v I__5116 (
            .O(N__21612),
            .I(N__21609));
    Span4Mux_h I__5115 (
            .O(N__21609),
            .I(N__21605));
    InMux I__5114 (
            .O(N__21608),
            .I(N__21602));
    Odrv4 I__5113 (
            .O(N__21605),
            .I(\Lab_UT.state_ret_11_RNI4RQC3_0 ));
    LocalMux I__5112 (
            .O(N__21602),
            .I(\Lab_UT.state_ret_11_RNI4RQC3_0 ));
    CascadeMux I__5111 (
            .O(N__21597),
            .I(\Lab_UT.state_ret_11_RNI4RQC3_0_cascade_ ));
    CascadeMux I__5110 (
            .O(N__21594),
            .I(N__21590));
    InMux I__5109 (
            .O(N__21593),
            .I(N__21585));
    InMux I__5108 (
            .O(N__21590),
            .I(N__21580));
    InMux I__5107 (
            .O(N__21589),
            .I(N__21580));
    IoInMux I__5106 (
            .O(N__21588),
            .I(N__21577));
    LocalMux I__5105 (
            .O(N__21585),
            .I(N__21574));
    LocalMux I__5104 (
            .O(N__21580),
            .I(N__21571));
    LocalMux I__5103 (
            .O(N__21577),
            .I(N__21567));
    Span4Mux_h I__5102 (
            .O(N__21574),
            .I(N__21562));
    Span4Mux_h I__5101 (
            .O(N__21571),
            .I(N__21562));
    InMux I__5100 (
            .O(N__21570),
            .I(N__21558));
    IoSpan4Mux I__5099 (
            .O(N__21567),
            .I(N__21555));
    Span4Mux_h I__5098 (
            .O(N__21562),
            .I(N__21552));
    InMux I__5097 (
            .O(N__21561),
            .I(N__21549));
    LocalMux I__5096 (
            .O(N__21558),
            .I(N__21546));
    Odrv4 I__5095 (
            .O(N__21555),
            .I(N_74));
    Odrv4 I__5094 (
            .O(N__21552),
            .I(N_74));
    LocalMux I__5093 (
            .O(N__21549),
            .I(N_74));
    Odrv4 I__5092 (
            .O(N__21546),
            .I(N_74));
    InMux I__5091 (
            .O(N__21537),
            .I(N__21531));
    InMux I__5090 (
            .O(N__21536),
            .I(N__21531));
    LocalMux I__5089 (
            .O(N__21531),
            .I(N__21528));
    Span4Mux_h I__5088 (
            .O(N__21528),
            .I(N__21525));
    Odrv4 I__5087 (
            .O(N__21525),
            .I(\Lab_UT.sccDnibble2En ));
    InMux I__5086 (
            .O(N__21522),
            .I(N__21515));
    InMux I__5085 (
            .O(N__21521),
            .I(N__21511));
    InMux I__5084 (
            .O(N__21520),
            .I(N__21508));
    InMux I__5083 (
            .O(N__21519),
            .I(N__21503));
    InMux I__5082 (
            .O(N__21518),
            .I(N__21503));
    LocalMux I__5081 (
            .O(N__21515),
            .I(N__21492));
    InMux I__5080 (
            .O(N__21514),
            .I(N__21489));
    LocalMux I__5079 (
            .O(N__21511),
            .I(N__21484));
    LocalMux I__5078 (
            .O(N__21508),
            .I(N__21484));
    LocalMux I__5077 (
            .O(N__21503),
            .I(N__21481));
    InMux I__5076 (
            .O(N__21502),
            .I(N__21472));
    InMux I__5075 (
            .O(N__21501),
            .I(N__21472));
    InMux I__5074 (
            .O(N__21500),
            .I(N__21472));
    InMux I__5073 (
            .O(N__21499),
            .I(N__21467));
    InMux I__5072 (
            .O(N__21498),
            .I(N__21467));
    InMux I__5071 (
            .O(N__21497),
            .I(N__21464));
    InMux I__5070 (
            .O(N__21496),
            .I(N__21459));
    InMux I__5069 (
            .O(N__21495),
            .I(N__21459));
    Span4Mux_h I__5068 (
            .O(N__21492),
            .I(N__21456));
    LocalMux I__5067 (
            .O(N__21489),
            .I(N__21453));
    Span4Mux_v I__5066 (
            .O(N__21484),
            .I(N__21448));
    Span4Mux_v I__5065 (
            .O(N__21481),
            .I(N__21448));
    InMux I__5064 (
            .O(N__21480),
            .I(N__21445));
    InMux I__5063 (
            .O(N__21479),
            .I(N__21442));
    LocalMux I__5062 (
            .O(N__21472),
            .I(N__21437));
    LocalMux I__5061 (
            .O(N__21467),
            .I(N__21437));
    LocalMux I__5060 (
            .O(N__21464),
            .I(N__21432));
    LocalMux I__5059 (
            .O(N__21459),
            .I(N__21432));
    Odrv4 I__5058 (
            .O(N__21456),
            .I(\Lab_UT.scctrl.N_223 ));
    Odrv4 I__5057 (
            .O(N__21453),
            .I(\Lab_UT.scctrl.N_223 ));
    Odrv4 I__5056 (
            .O(N__21448),
            .I(\Lab_UT.scctrl.N_223 ));
    LocalMux I__5055 (
            .O(N__21445),
            .I(\Lab_UT.scctrl.N_223 ));
    LocalMux I__5054 (
            .O(N__21442),
            .I(\Lab_UT.scctrl.N_223 ));
    Odrv4 I__5053 (
            .O(N__21437),
            .I(\Lab_UT.scctrl.N_223 ));
    Odrv12 I__5052 (
            .O(N__21432),
            .I(\Lab_UT.scctrl.N_223 ));
    CascadeMux I__5051 (
            .O(N__21417),
            .I(N__21405));
    InMux I__5050 (
            .O(N__21416),
            .I(N__21399));
    InMux I__5049 (
            .O(N__21415),
            .I(N__21392));
    InMux I__5048 (
            .O(N__21414),
            .I(N__21392));
    InMux I__5047 (
            .O(N__21413),
            .I(N__21392));
    InMux I__5046 (
            .O(N__21412),
            .I(N__21381));
    InMux I__5045 (
            .O(N__21411),
            .I(N__21381));
    InMux I__5044 (
            .O(N__21410),
            .I(N__21381));
    CascadeMux I__5043 (
            .O(N__21409),
            .I(N__21378));
    InMux I__5042 (
            .O(N__21408),
            .I(N__21374));
    InMux I__5041 (
            .O(N__21405),
            .I(N__21371));
    InMux I__5040 (
            .O(N__21404),
            .I(N__21366));
    InMux I__5039 (
            .O(N__21403),
            .I(N__21359));
    InMux I__5038 (
            .O(N__21402),
            .I(N__21359));
    LocalMux I__5037 (
            .O(N__21399),
            .I(N__21356));
    LocalMux I__5036 (
            .O(N__21392),
            .I(N__21353));
    InMux I__5035 (
            .O(N__21391),
            .I(N__21350));
    InMux I__5034 (
            .O(N__21390),
            .I(N__21347));
    InMux I__5033 (
            .O(N__21389),
            .I(N__21342));
    InMux I__5032 (
            .O(N__21388),
            .I(N__21342));
    LocalMux I__5031 (
            .O(N__21381),
            .I(N__21339));
    InMux I__5030 (
            .O(N__21378),
            .I(N__21334));
    InMux I__5029 (
            .O(N__21377),
            .I(N__21334));
    LocalMux I__5028 (
            .O(N__21374),
            .I(N__21329));
    LocalMux I__5027 (
            .O(N__21371),
            .I(N__21326));
    InMux I__5026 (
            .O(N__21370),
            .I(N__21321));
    InMux I__5025 (
            .O(N__21369),
            .I(N__21321));
    LocalMux I__5024 (
            .O(N__21366),
            .I(N__21318));
    InMux I__5023 (
            .O(N__21365),
            .I(N__21309));
    InMux I__5022 (
            .O(N__21364),
            .I(N__21309));
    LocalMux I__5021 (
            .O(N__21359),
            .I(N__21306));
    Span4Mux_v I__5020 (
            .O(N__21356),
            .I(N__21300));
    Span4Mux_v I__5019 (
            .O(N__21353),
            .I(N__21300));
    LocalMux I__5018 (
            .O(N__21350),
            .I(N__21297));
    LocalMux I__5017 (
            .O(N__21347),
            .I(N__21288));
    LocalMux I__5016 (
            .O(N__21342),
            .I(N__21288));
    Span4Mux_v I__5015 (
            .O(N__21339),
            .I(N__21288));
    LocalMux I__5014 (
            .O(N__21334),
            .I(N__21288));
    InMux I__5013 (
            .O(N__21333),
            .I(N__21283));
    InMux I__5012 (
            .O(N__21332),
            .I(N__21283));
    Span4Mux_v I__5011 (
            .O(N__21329),
            .I(N__21280));
    Span4Mux_v I__5010 (
            .O(N__21326),
            .I(N__21275));
    LocalMux I__5009 (
            .O(N__21321),
            .I(N__21275));
    Span4Mux_s2_h I__5008 (
            .O(N__21318),
            .I(N__21272));
    InMux I__5007 (
            .O(N__21317),
            .I(N__21267));
    InMux I__5006 (
            .O(N__21316),
            .I(N__21267));
    InMux I__5005 (
            .O(N__21315),
            .I(N__21264));
    InMux I__5004 (
            .O(N__21314),
            .I(N__21261));
    LocalMux I__5003 (
            .O(N__21309),
            .I(N__21258));
    Span4Mux_s3_h I__5002 (
            .O(N__21306),
            .I(N__21255));
    InMux I__5001 (
            .O(N__21305),
            .I(N__21252));
    Span4Mux_h I__5000 (
            .O(N__21300),
            .I(N__21243));
    Span4Mux_h I__4999 (
            .O(N__21297),
            .I(N__21243));
    Span4Mux_v I__4998 (
            .O(N__21288),
            .I(N__21243));
    LocalMux I__4997 (
            .O(N__21283),
            .I(N__21243));
    Span4Mux_v I__4996 (
            .O(N__21280),
            .I(N__21236));
    Span4Mux_v I__4995 (
            .O(N__21275),
            .I(N__21236));
    Span4Mux_v I__4994 (
            .O(N__21272),
            .I(N__21236));
    LocalMux I__4993 (
            .O(N__21267),
            .I(\Lab_UT.scctrl.stateZ0Z_0 ));
    LocalMux I__4992 (
            .O(N__21264),
            .I(\Lab_UT.scctrl.stateZ0Z_0 ));
    LocalMux I__4991 (
            .O(N__21261),
            .I(\Lab_UT.scctrl.stateZ0Z_0 ));
    Odrv4 I__4990 (
            .O(N__21258),
            .I(\Lab_UT.scctrl.stateZ0Z_0 ));
    Odrv4 I__4989 (
            .O(N__21255),
            .I(\Lab_UT.scctrl.stateZ0Z_0 ));
    LocalMux I__4988 (
            .O(N__21252),
            .I(\Lab_UT.scctrl.stateZ0Z_0 ));
    Odrv4 I__4987 (
            .O(N__21243),
            .I(\Lab_UT.scctrl.stateZ0Z_0 ));
    Odrv4 I__4986 (
            .O(N__21236),
            .I(\Lab_UT.scctrl.stateZ0Z_0 ));
    CascadeMux I__4985 (
            .O(N__21219),
            .I(N__21216));
    InMux I__4984 (
            .O(N__21216),
            .I(N__21213));
    LocalMux I__4983 (
            .O(N__21213),
            .I(N__21210));
    Span4Mux_v I__4982 (
            .O(N__21210),
            .I(N__21207));
    Odrv4 I__4981 (
            .O(N__21207),
            .I(\Lab_UT.scctrl.N_5_0 ));
    InMux I__4980 (
            .O(N__21204),
            .I(N__21201));
    LocalMux I__4979 (
            .O(N__21201),
            .I(N__21198));
    Span4Mux_v I__4978 (
            .O(N__21198),
            .I(N__21195));
    Odrv4 I__4977 (
            .O(N__21195),
            .I(\Lab_UT.scctrl.G_10_i_a7_0_2 ));
    IoInMux I__4976 (
            .O(N__21192),
            .I(N__21189));
    LocalMux I__4975 (
            .O(N__21189),
            .I(N__21184));
    InMux I__4974 (
            .O(N__21188),
            .I(N__21181));
    InMux I__4973 (
            .O(N__21187),
            .I(N__21178));
    Span4Mux_s1_v I__4972 (
            .O(N__21184),
            .I(N__21175));
    LocalMux I__4971 (
            .O(N__21181),
            .I(N__21172));
    LocalMux I__4970 (
            .O(N__21178),
            .I(N__21169));
    Span4Mux_v I__4969 (
            .O(N__21175),
            .I(N__21166));
    Span4Mux_v I__4968 (
            .O(N__21172),
            .I(N__21161));
    Span4Mux_s1_h I__4967 (
            .O(N__21169),
            .I(N__21161));
    Span4Mux_h I__4966 (
            .O(N__21166),
            .I(N__21158));
    Span4Mux_h I__4965 (
            .O(N__21161),
            .I(N__21155));
    Odrv4 I__4964 (
            .O(N__21158),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4963 (
            .O(N__21155),
            .I(CONSTANT_ONE_NET));
    ClkMux I__4962 (
            .O(N__21150),
            .I(N__20907));
    ClkMux I__4961 (
            .O(N__21149),
            .I(N__20907));
    ClkMux I__4960 (
            .O(N__21148),
            .I(N__20907));
    ClkMux I__4959 (
            .O(N__21147),
            .I(N__20907));
    ClkMux I__4958 (
            .O(N__21146),
            .I(N__20907));
    ClkMux I__4957 (
            .O(N__21145),
            .I(N__20907));
    ClkMux I__4956 (
            .O(N__21144),
            .I(N__20907));
    ClkMux I__4955 (
            .O(N__21143),
            .I(N__20907));
    ClkMux I__4954 (
            .O(N__21142),
            .I(N__20907));
    ClkMux I__4953 (
            .O(N__21141),
            .I(N__20907));
    ClkMux I__4952 (
            .O(N__21140),
            .I(N__20907));
    ClkMux I__4951 (
            .O(N__21139),
            .I(N__20907));
    ClkMux I__4950 (
            .O(N__21138),
            .I(N__20907));
    ClkMux I__4949 (
            .O(N__21137),
            .I(N__20907));
    ClkMux I__4948 (
            .O(N__21136),
            .I(N__20907));
    ClkMux I__4947 (
            .O(N__21135),
            .I(N__20907));
    ClkMux I__4946 (
            .O(N__21134),
            .I(N__20907));
    ClkMux I__4945 (
            .O(N__21133),
            .I(N__20907));
    ClkMux I__4944 (
            .O(N__21132),
            .I(N__20907));
    ClkMux I__4943 (
            .O(N__21131),
            .I(N__20907));
    ClkMux I__4942 (
            .O(N__21130),
            .I(N__20907));
    ClkMux I__4941 (
            .O(N__21129),
            .I(N__20907));
    ClkMux I__4940 (
            .O(N__21128),
            .I(N__20907));
    ClkMux I__4939 (
            .O(N__21127),
            .I(N__20907));
    ClkMux I__4938 (
            .O(N__21126),
            .I(N__20907));
    ClkMux I__4937 (
            .O(N__21125),
            .I(N__20907));
    ClkMux I__4936 (
            .O(N__21124),
            .I(N__20907));
    ClkMux I__4935 (
            .O(N__21123),
            .I(N__20907));
    ClkMux I__4934 (
            .O(N__21122),
            .I(N__20907));
    ClkMux I__4933 (
            .O(N__21121),
            .I(N__20907));
    ClkMux I__4932 (
            .O(N__21120),
            .I(N__20907));
    ClkMux I__4931 (
            .O(N__21119),
            .I(N__20907));
    ClkMux I__4930 (
            .O(N__21118),
            .I(N__20907));
    ClkMux I__4929 (
            .O(N__21117),
            .I(N__20907));
    ClkMux I__4928 (
            .O(N__21116),
            .I(N__20907));
    ClkMux I__4927 (
            .O(N__21115),
            .I(N__20907));
    ClkMux I__4926 (
            .O(N__21114),
            .I(N__20907));
    ClkMux I__4925 (
            .O(N__21113),
            .I(N__20907));
    ClkMux I__4924 (
            .O(N__21112),
            .I(N__20907));
    ClkMux I__4923 (
            .O(N__21111),
            .I(N__20907));
    ClkMux I__4922 (
            .O(N__21110),
            .I(N__20907));
    ClkMux I__4921 (
            .O(N__21109),
            .I(N__20907));
    ClkMux I__4920 (
            .O(N__21108),
            .I(N__20907));
    ClkMux I__4919 (
            .O(N__21107),
            .I(N__20907));
    ClkMux I__4918 (
            .O(N__21106),
            .I(N__20907));
    ClkMux I__4917 (
            .O(N__21105),
            .I(N__20907));
    ClkMux I__4916 (
            .O(N__21104),
            .I(N__20907));
    ClkMux I__4915 (
            .O(N__21103),
            .I(N__20907));
    ClkMux I__4914 (
            .O(N__21102),
            .I(N__20907));
    ClkMux I__4913 (
            .O(N__21101),
            .I(N__20907));
    ClkMux I__4912 (
            .O(N__21100),
            .I(N__20907));
    ClkMux I__4911 (
            .O(N__21099),
            .I(N__20907));
    ClkMux I__4910 (
            .O(N__21098),
            .I(N__20907));
    ClkMux I__4909 (
            .O(N__21097),
            .I(N__20907));
    ClkMux I__4908 (
            .O(N__21096),
            .I(N__20907));
    ClkMux I__4907 (
            .O(N__21095),
            .I(N__20907));
    ClkMux I__4906 (
            .O(N__21094),
            .I(N__20907));
    ClkMux I__4905 (
            .O(N__21093),
            .I(N__20907));
    ClkMux I__4904 (
            .O(N__21092),
            .I(N__20907));
    ClkMux I__4903 (
            .O(N__21091),
            .I(N__20907));
    ClkMux I__4902 (
            .O(N__21090),
            .I(N__20907));
    ClkMux I__4901 (
            .O(N__21089),
            .I(N__20907));
    ClkMux I__4900 (
            .O(N__21088),
            .I(N__20907));
    ClkMux I__4899 (
            .O(N__21087),
            .I(N__20907));
    ClkMux I__4898 (
            .O(N__21086),
            .I(N__20907));
    ClkMux I__4897 (
            .O(N__21085),
            .I(N__20907));
    ClkMux I__4896 (
            .O(N__21084),
            .I(N__20907));
    ClkMux I__4895 (
            .O(N__21083),
            .I(N__20907));
    ClkMux I__4894 (
            .O(N__21082),
            .I(N__20907));
    ClkMux I__4893 (
            .O(N__21081),
            .I(N__20907));
    ClkMux I__4892 (
            .O(N__21080),
            .I(N__20907));
    ClkMux I__4891 (
            .O(N__21079),
            .I(N__20907));
    ClkMux I__4890 (
            .O(N__21078),
            .I(N__20907));
    ClkMux I__4889 (
            .O(N__21077),
            .I(N__20907));
    ClkMux I__4888 (
            .O(N__21076),
            .I(N__20907));
    ClkMux I__4887 (
            .O(N__21075),
            .I(N__20907));
    ClkMux I__4886 (
            .O(N__21074),
            .I(N__20907));
    ClkMux I__4885 (
            .O(N__21073),
            .I(N__20907));
    ClkMux I__4884 (
            .O(N__21072),
            .I(N__20907));
    ClkMux I__4883 (
            .O(N__21071),
            .I(N__20907));
    ClkMux I__4882 (
            .O(N__21070),
            .I(N__20907));
    GlobalMux I__4881 (
            .O(N__20907),
            .I(N__20904));
    gio2CtrlBuf I__4880 (
            .O(N__20904),
            .I(clk_g));
    CEMux I__4879 (
            .O(N__20901),
            .I(N__20896));
    CEMux I__4878 (
            .O(N__20900),
            .I(N__20893));
    CEMux I__4877 (
            .O(N__20899),
            .I(N__20889));
    LocalMux I__4876 (
            .O(N__20896),
            .I(N__20886));
    LocalMux I__4875 (
            .O(N__20893),
            .I(N__20883));
    CEMux I__4874 (
            .O(N__20892),
            .I(N__20880));
    LocalMux I__4873 (
            .O(N__20889),
            .I(N__20877));
    Span4Mux_h I__4872 (
            .O(N__20886),
            .I(N__20874));
    Span4Mux_h I__4871 (
            .O(N__20883),
            .I(N__20869));
    LocalMux I__4870 (
            .O(N__20880),
            .I(N__20869));
    Odrv4 I__4869 (
            .O(N__20877),
            .I(\Lab_UT.scctrl.next_state_RNIN96CP1Z0Z_3 ));
    Odrv4 I__4868 (
            .O(N__20874),
            .I(\Lab_UT.scctrl.next_state_RNIN96CP1Z0Z_3 ));
    Odrv4 I__4867 (
            .O(N__20869),
            .I(\Lab_UT.scctrl.next_state_RNIN96CP1Z0Z_3 ));
    InMux I__4866 (
            .O(N__20862),
            .I(N__20859));
    LocalMux I__4865 (
            .O(N__20859),
            .I(N__20804));
    SRMux I__4864 (
            .O(N__20858),
            .I(N__20697));
    SRMux I__4863 (
            .O(N__20857),
            .I(N__20697));
    SRMux I__4862 (
            .O(N__20856),
            .I(N__20697));
    SRMux I__4861 (
            .O(N__20855),
            .I(N__20697));
    SRMux I__4860 (
            .O(N__20854),
            .I(N__20697));
    SRMux I__4859 (
            .O(N__20853),
            .I(N__20697));
    SRMux I__4858 (
            .O(N__20852),
            .I(N__20697));
    SRMux I__4857 (
            .O(N__20851),
            .I(N__20697));
    SRMux I__4856 (
            .O(N__20850),
            .I(N__20697));
    SRMux I__4855 (
            .O(N__20849),
            .I(N__20697));
    SRMux I__4854 (
            .O(N__20848),
            .I(N__20697));
    SRMux I__4853 (
            .O(N__20847),
            .I(N__20697));
    SRMux I__4852 (
            .O(N__20846),
            .I(N__20697));
    SRMux I__4851 (
            .O(N__20845),
            .I(N__20697));
    SRMux I__4850 (
            .O(N__20844),
            .I(N__20697));
    SRMux I__4849 (
            .O(N__20843),
            .I(N__20697));
    SRMux I__4848 (
            .O(N__20842),
            .I(N__20697));
    SRMux I__4847 (
            .O(N__20841),
            .I(N__20697));
    SRMux I__4846 (
            .O(N__20840),
            .I(N__20697));
    SRMux I__4845 (
            .O(N__20839),
            .I(N__20697));
    SRMux I__4844 (
            .O(N__20838),
            .I(N__20697));
    SRMux I__4843 (
            .O(N__20837),
            .I(N__20697));
    SRMux I__4842 (
            .O(N__20836),
            .I(N__20697));
    SRMux I__4841 (
            .O(N__20835),
            .I(N__20697));
    SRMux I__4840 (
            .O(N__20834),
            .I(N__20697));
    SRMux I__4839 (
            .O(N__20833),
            .I(N__20697));
    SRMux I__4838 (
            .O(N__20832),
            .I(N__20697));
    SRMux I__4837 (
            .O(N__20831),
            .I(N__20697));
    SRMux I__4836 (
            .O(N__20830),
            .I(N__20697));
    SRMux I__4835 (
            .O(N__20829),
            .I(N__20697));
    SRMux I__4834 (
            .O(N__20828),
            .I(N__20697));
    SRMux I__4833 (
            .O(N__20827),
            .I(N__20697));
    SRMux I__4832 (
            .O(N__20826),
            .I(N__20697));
    SRMux I__4831 (
            .O(N__20825),
            .I(N__20697));
    SRMux I__4830 (
            .O(N__20824),
            .I(N__20697));
    SRMux I__4829 (
            .O(N__20823),
            .I(N__20697));
    SRMux I__4828 (
            .O(N__20822),
            .I(N__20697));
    SRMux I__4827 (
            .O(N__20821),
            .I(N__20697));
    SRMux I__4826 (
            .O(N__20820),
            .I(N__20697));
    SRMux I__4825 (
            .O(N__20819),
            .I(N__20697));
    SRMux I__4824 (
            .O(N__20818),
            .I(N__20697));
    SRMux I__4823 (
            .O(N__20817),
            .I(N__20697));
    SRMux I__4822 (
            .O(N__20816),
            .I(N__20697));
    SRMux I__4821 (
            .O(N__20815),
            .I(N__20697));
    SRMux I__4820 (
            .O(N__20814),
            .I(N__20697));
    SRMux I__4819 (
            .O(N__20813),
            .I(N__20697));
    SRMux I__4818 (
            .O(N__20812),
            .I(N__20697));
    SRMux I__4817 (
            .O(N__20811),
            .I(N__20697));
    SRMux I__4816 (
            .O(N__20810),
            .I(N__20697));
    SRMux I__4815 (
            .O(N__20809),
            .I(N__20697));
    SRMux I__4814 (
            .O(N__20808),
            .I(N__20697));
    SRMux I__4813 (
            .O(N__20807),
            .I(N__20697));
    Glb2LocalMux I__4812 (
            .O(N__20804),
            .I(N__20697));
    GlobalMux I__4811 (
            .O(N__20697),
            .I(N__20694));
    gio2CtrlBuf I__4810 (
            .O(N__20694),
            .I(resetGen_rst_1_iso_g));
    CascadeMux I__4809 (
            .O(N__20691),
            .I(N__20687));
    InMux I__4808 (
            .O(N__20690),
            .I(N__20681));
    InMux I__4807 (
            .O(N__20687),
            .I(N__20681));
    InMux I__4806 (
            .O(N__20686),
            .I(N__20678));
    LocalMux I__4805 (
            .O(N__20681),
            .I(N__20675));
    LocalMux I__4804 (
            .O(N__20678),
            .I(N__20672));
    Span4Mux_v I__4803 (
            .O(N__20675),
            .I(N__20669));
    Odrv4 I__4802 (
            .O(N__20672),
            .I(\Lab_UT.scctrl.N_260 ));
    Odrv4 I__4801 (
            .O(N__20669),
            .I(\Lab_UT.scctrl.N_260 ));
    InMux I__4800 (
            .O(N__20664),
            .I(N__20658));
    InMux I__4799 (
            .O(N__20663),
            .I(N__20652));
    CascadeMux I__4798 (
            .O(N__20662),
            .I(N__20648));
    CascadeMux I__4797 (
            .O(N__20661),
            .I(N__20644));
    LocalMux I__4796 (
            .O(N__20658),
            .I(N__20638));
    InMux I__4795 (
            .O(N__20657),
            .I(N__20635));
    InMux I__4794 (
            .O(N__20656),
            .I(N__20632));
    InMux I__4793 (
            .O(N__20655),
            .I(N__20629));
    LocalMux I__4792 (
            .O(N__20652),
            .I(N__20626));
    InMux I__4791 (
            .O(N__20651),
            .I(N__20623));
    InMux I__4790 (
            .O(N__20648),
            .I(N__20620));
    InMux I__4789 (
            .O(N__20647),
            .I(N__20617));
    InMux I__4788 (
            .O(N__20644),
            .I(N__20614));
    InMux I__4787 (
            .O(N__20643),
            .I(N__20609));
    InMux I__4786 (
            .O(N__20642),
            .I(N__20609));
    InMux I__4785 (
            .O(N__20641),
            .I(N__20606));
    Span4Mux_h I__4784 (
            .O(N__20638),
            .I(N__20596));
    LocalMux I__4783 (
            .O(N__20635),
            .I(N__20596));
    LocalMux I__4782 (
            .O(N__20632),
            .I(N__20596));
    LocalMux I__4781 (
            .O(N__20629),
            .I(N__20596));
    Span4Mux_h I__4780 (
            .O(N__20626),
            .I(N__20591));
    LocalMux I__4779 (
            .O(N__20623),
            .I(N__20591));
    LocalMux I__4778 (
            .O(N__20620),
            .I(N__20586));
    LocalMux I__4777 (
            .O(N__20617),
            .I(N__20586));
    LocalMux I__4776 (
            .O(N__20614),
            .I(N__20578));
    LocalMux I__4775 (
            .O(N__20609),
            .I(N__20578));
    LocalMux I__4774 (
            .O(N__20606),
            .I(N__20578));
    CascadeMux I__4773 (
            .O(N__20605),
            .I(N__20574));
    Sp12to4 I__4772 (
            .O(N__20596),
            .I(N__20571));
    Span4Mux_v I__4771 (
            .O(N__20591),
            .I(N__20566));
    Span4Mux_v I__4770 (
            .O(N__20586),
            .I(N__20566));
    InMux I__4769 (
            .O(N__20585),
            .I(N__20563));
    Span4Mux_h I__4768 (
            .O(N__20578),
            .I(N__20560));
    InMux I__4767 (
            .O(N__20577),
            .I(N__20557));
    InMux I__4766 (
            .O(N__20574),
            .I(N__20554));
    Odrv12 I__4765 (
            .O(N__20571),
            .I(\Lab_UT.scctrl.N_235 ));
    Odrv4 I__4764 (
            .O(N__20566),
            .I(\Lab_UT.scctrl.N_235 ));
    LocalMux I__4763 (
            .O(N__20563),
            .I(\Lab_UT.scctrl.N_235 ));
    Odrv4 I__4762 (
            .O(N__20560),
            .I(\Lab_UT.scctrl.N_235 ));
    LocalMux I__4761 (
            .O(N__20557),
            .I(\Lab_UT.scctrl.N_235 ));
    LocalMux I__4760 (
            .O(N__20554),
            .I(\Lab_UT.scctrl.N_235 ));
    IoInMux I__4759 (
            .O(N__20541),
            .I(N__20538));
    LocalMux I__4758 (
            .O(N__20538),
            .I(N__20535));
    IoSpan4Mux I__4757 (
            .O(N__20535),
            .I(N__20532));
    Odrv4 I__4756 (
            .O(N__20532),
            .I(N_55_i));
    CascadeMux I__4755 (
            .O(N__20529),
            .I(N__20525));
    InMux I__4754 (
            .O(N__20528),
            .I(N__20517));
    InMux I__4753 (
            .O(N__20525),
            .I(N__20514));
    InMux I__4752 (
            .O(N__20524),
            .I(N__20509));
    InMux I__4751 (
            .O(N__20523),
            .I(N__20505));
    InMux I__4750 (
            .O(N__20522),
            .I(N__20502));
    InMux I__4749 (
            .O(N__20521),
            .I(N__20499));
    InMux I__4748 (
            .O(N__20520),
            .I(N__20496));
    LocalMux I__4747 (
            .O(N__20517),
            .I(N__20491));
    LocalMux I__4746 (
            .O(N__20514),
            .I(N__20491));
    InMux I__4745 (
            .O(N__20513),
            .I(N__20486));
    InMux I__4744 (
            .O(N__20512),
            .I(N__20486));
    LocalMux I__4743 (
            .O(N__20509),
            .I(N__20483));
    InMux I__4742 (
            .O(N__20508),
            .I(N__20480));
    LocalMux I__4741 (
            .O(N__20505),
            .I(N__20475));
    LocalMux I__4740 (
            .O(N__20502),
            .I(N__20475));
    LocalMux I__4739 (
            .O(N__20499),
            .I(N__20472));
    LocalMux I__4738 (
            .O(N__20496),
            .I(\Lab_UT.scctrl.state_i_1_0_rep1 ));
    Odrv4 I__4737 (
            .O(N__20491),
            .I(\Lab_UT.scctrl.state_i_1_0_rep1 ));
    LocalMux I__4736 (
            .O(N__20486),
            .I(\Lab_UT.scctrl.state_i_1_0_rep1 ));
    Odrv12 I__4735 (
            .O(N__20483),
            .I(\Lab_UT.scctrl.state_i_1_0_rep1 ));
    LocalMux I__4734 (
            .O(N__20480),
            .I(\Lab_UT.scctrl.state_i_1_0_rep1 ));
    Odrv4 I__4733 (
            .O(N__20475),
            .I(\Lab_UT.scctrl.state_i_1_0_rep1 ));
    Odrv4 I__4732 (
            .O(N__20472),
            .I(\Lab_UT.scctrl.state_i_1_0_rep1 ));
    CascadeMux I__4731 (
            .O(N__20457),
            .I(N__20453));
    CascadeMux I__4730 (
            .O(N__20456),
            .I(N__20448));
    InMux I__4729 (
            .O(N__20453),
            .I(N__20444));
    InMux I__4728 (
            .O(N__20452),
            .I(N__20441));
    InMux I__4727 (
            .O(N__20451),
            .I(N__20438));
    InMux I__4726 (
            .O(N__20448),
            .I(N__20435));
    CascadeMux I__4725 (
            .O(N__20447),
            .I(N__20430));
    LocalMux I__4724 (
            .O(N__20444),
            .I(N__20427));
    LocalMux I__4723 (
            .O(N__20441),
            .I(N__20424));
    LocalMux I__4722 (
            .O(N__20438),
            .I(N__20419));
    LocalMux I__4721 (
            .O(N__20435),
            .I(N__20419));
    InMux I__4720 (
            .O(N__20434),
            .I(N__20414));
    InMux I__4719 (
            .O(N__20433),
            .I(N__20414));
    InMux I__4718 (
            .O(N__20430),
            .I(N__20411));
    Span4Mux_h I__4717 (
            .O(N__20427),
            .I(N__20404));
    Span4Mux_h I__4716 (
            .O(N__20424),
            .I(N__20404));
    Span4Mux_v I__4715 (
            .O(N__20419),
            .I(N__20404));
    LocalMux I__4714 (
            .O(N__20414),
            .I(N__20399));
    LocalMux I__4713 (
            .O(N__20411),
            .I(N__20399));
    Span4Mux_v I__4712 (
            .O(N__20404),
            .I(N__20394));
    Span4Mux_v I__4711 (
            .O(N__20399),
            .I(N__20394));
    Odrv4 I__4710 (
            .O(N__20394),
            .I(\Lab_UT.scctrl.state_2_rep1 ));
    InMux I__4709 (
            .O(N__20391),
            .I(N__20388));
    LocalMux I__4708 (
            .O(N__20388),
            .I(\Lab_UT.scctrl.N_13_1 ));
    CascadeMux I__4707 (
            .O(N__20385),
            .I(\Lab_UT.scctrl.G_10_i_1_cascade_ ));
    InMux I__4706 (
            .O(N__20382),
            .I(N__20379));
    LocalMux I__4705 (
            .O(N__20379),
            .I(N__20376));
    Span4Mux_s2_h I__4704 (
            .O(N__20376),
            .I(N__20372));
    InMux I__4703 (
            .O(N__20375),
            .I(N__20369));
    Span4Mux_v I__4702 (
            .O(N__20372),
            .I(N__20366));
    LocalMux I__4701 (
            .O(N__20369),
            .I(N__20363));
    Odrv4 I__4700 (
            .O(N__20366),
            .I(\Lab_UT.scctrl.state_fast_2 ));
    Odrv12 I__4699 (
            .O(N__20363),
            .I(\Lab_UT.scctrl.state_fast_2 ));
    InMux I__4698 (
            .O(N__20358),
            .I(N__20355));
    LocalMux I__4697 (
            .O(N__20355),
            .I(N__20351));
    InMux I__4696 (
            .O(N__20354),
            .I(N__20347));
    Span4Mux_s3_h I__4695 (
            .O(N__20351),
            .I(N__20344));
    InMux I__4694 (
            .O(N__20350),
            .I(N__20341));
    LocalMux I__4693 (
            .O(N__20347),
            .I(N__20338));
    Odrv4 I__4692 (
            .O(N__20344),
            .I(\Lab_UT.scctrl.state_i_1_fast_0 ));
    LocalMux I__4691 (
            .O(N__20341),
            .I(\Lab_UT.scctrl.state_i_1_fast_0 ));
    Odrv12 I__4690 (
            .O(N__20338),
            .I(\Lab_UT.scctrl.state_i_1_fast_0 ));
    CascadeMux I__4689 (
            .O(N__20331),
            .I(\Lab_UT.scctrl.next_state_1_0_cascade_ ));
    CascadeMux I__4688 (
            .O(N__20328),
            .I(N__20325));
    InMux I__4687 (
            .O(N__20325),
            .I(N__20322));
    LocalMux I__4686 (
            .O(N__20322),
            .I(N__20319));
    Span4Mux_h I__4685 (
            .O(N__20319),
            .I(N__20316));
    Odrv4 I__4684 (
            .O(N__20316),
            .I(\Lab_UT.scctrl.N_356_1_0 ));
    InMux I__4683 (
            .O(N__20313),
            .I(N__20310));
    LocalMux I__4682 (
            .O(N__20310),
            .I(N__20307));
    Span4Mux_h I__4681 (
            .O(N__20307),
            .I(N__20304));
    Odrv4 I__4680 (
            .O(N__20304),
            .I(\Lab_UT.scctrl.g0_9_a2_1 ));
    InMux I__4679 (
            .O(N__20301),
            .I(N__20298));
    LocalMux I__4678 (
            .O(N__20298),
            .I(N__20295));
    Span4Mux_s3_h I__4677 (
            .O(N__20295),
            .I(N__20292));
    Odrv4 I__4676 (
            .O(N__20292),
            .I(\Lab_UT.scctrl.g0_2_3_1 ));
    CascadeMux I__4675 (
            .O(N__20289),
            .I(N__20280));
    CascadeMux I__4674 (
            .O(N__20288),
            .I(N__20277));
    CascadeMux I__4673 (
            .O(N__20287),
            .I(N__20273));
    CascadeMux I__4672 (
            .O(N__20286),
            .I(N__20270));
    InMux I__4671 (
            .O(N__20285),
            .I(N__20262));
    InMux I__4670 (
            .O(N__20284),
            .I(N__20262));
    CascadeMux I__4669 (
            .O(N__20283),
            .I(N__20259));
    InMux I__4668 (
            .O(N__20280),
            .I(N__20253));
    InMux I__4667 (
            .O(N__20277),
            .I(N__20253));
    InMux I__4666 (
            .O(N__20276),
            .I(N__20247));
    InMux I__4665 (
            .O(N__20273),
            .I(N__20236));
    InMux I__4664 (
            .O(N__20270),
            .I(N__20236));
    InMux I__4663 (
            .O(N__20269),
            .I(N__20236));
    InMux I__4662 (
            .O(N__20268),
            .I(N__20236));
    InMux I__4661 (
            .O(N__20267),
            .I(N__20236));
    LocalMux I__4660 (
            .O(N__20262),
            .I(N__20233));
    InMux I__4659 (
            .O(N__20259),
            .I(N__20228));
    InMux I__4658 (
            .O(N__20258),
            .I(N__20228));
    LocalMux I__4657 (
            .O(N__20253),
            .I(N__20225));
    InMux I__4656 (
            .O(N__20252),
            .I(N__20218));
    InMux I__4655 (
            .O(N__20251),
            .I(N__20218));
    InMux I__4654 (
            .O(N__20250),
            .I(N__20218));
    LocalMux I__4653 (
            .O(N__20247),
            .I(N__20209));
    LocalMux I__4652 (
            .O(N__20236),
            .I(N__20209));
    Span4Mux_v I__4651 (
            .O(N__20233),
            .I(N__20209));
    LocalMux I__4650 (
            .O(N__20228),
            .I(N__20209));
    Span4Mux_v I__4649 (
            .O(N__20225),
            .I(N__20204));
    LocalMux I__4648 (
            .O(N__20218),
            .I(N__20204));
    Span4Mux_v I__4647 (
            .O(N__20209),
            .I(N__20199));
    Span4Mux_h I__4646 (
            .O(N__20204),
            .I(N__20199));
    Odrv4 I__4645 (
            .O(N__20199),
            .I(\Lab_UT.scctrl.next_stateZ0Z_0 ));
    InMux I__4644 (
            .O(N__20196),
            .I(N__20193));
    LocalMux I__4643 (
            .O(N__20193),
            .I(N__20190));
    Span4Mux_h I__4642 (
            .O(N__20190),
            .I(N__20187));
    Odrv4 I__4641 (
            .O(N__20187),
            .I(\Lab_UT.scctrl.g0_2_2_1 ));
    InMux I__4640 (
            .O(N__20184),
            .I(N__20172));
    InMux I__4639 (
            .O(N__20183),
            .I(N__20169));
    InMux I__4638 (
            .O(N__20182),
            .I(N__20166));
    InMux I__4637 (
            .O(N__20181),
            .I(N__20161));
    InMux I__4636 (
            .O(N__20180),
            .I(N__20161));
    InMux I__4635 (
            .O(N__20179),
            .I(N__20158));
    InMux I__4634 (
            .O(N__20178),
            .I(N__20151));
    InMux I__4633 (
            .O(N__20177),
            .I(N__20151));
    InMux I__4632 (
            .O(N__20176),
            .I(N__20151));
    InMux I__4631 (
            .O(N__20175),
            .I(N__20148));
    LocalMux I__4630 (
            .O(N__20172),
            .I(N__20145));
    LocalMux I__4629 (
            .O(N__20169),
            .I(N__20142));
    LocalMux I__4628 (
            .O(N__20166),
            .I(N__20136));
    LocalMux I__4627 (
            .O(N__20161),
            .I(N__20131));
    LocalMux I__4626 (
            .O(N__20158),
            .I(N__20131));
    LocalMux I__4625 (
            .O(N__20151),
            .I(N__20128));
    LocalMux I__4624 (
            .O(N__20148),
            .I(N__20125));
    Span4Mux_v I__4623 (
            .O(N__20145),
            .I(N__20122));
    Span4Mux_h I__4622 (
            .O(N__20142),
            .I(N__20119));
    CascadeMux I__4621 (
            .O(N__20141),
            .I(N__20115));
    InMux I__4620 (
            .O(N__20140),
            .I(N__20111));
    InMux I__4619 (
            .O(N__20139),
            .I(N__20108));
    Span4Mux_v I__4618 (
            .O(N__20136),
            .I(N__20103));
    Span4Mux_v I__4617 (
            .O(N__20131),
            .I(N__20103));
    Span4Mux_h I__4616 (
            .O(N__20128),
            .I(N__20100));
    Span4Mux_v I__4615 (
            .O(N__20125),
            .I(N__20097));
    Span4Mux_h I__4614 (
            .O(N__20122),
            .I(N__20092));
    Span4Mux_v I__4613 (
            .O(N__20119),
            .I(N__20092));
    InMux I__4612 (
            .O(N__20118),
            .I(N__20089));
    InMux I__4611 (
            .O(N__20115),
            .I(N__20084));
    InMux I__4610 (
            .O(N__20114),
            .I(N__20084));
    LocalMux I__4609 (
            .O(N__20111),
            .I(N__20079));
    LocalMux I__4608 (
            .O(N__20108),
            .I(N__20079));
    Span4Mux_h I__4607 (
            .O(N__20103),
            .I(N__20076));
    Odrv4 I__4606 (
            .O(N__20100),
            .I(rst));
    Odrv4 I__4605 (
            .O(N__20097),
            .I(rst));
    Odrv4 I__4604 (
            .O(N__20092),
            .I(rst));
    LocalMux I__4603 (
            .O(N__20089),
            .I(rst));
    LocalMux I__4602 (
            .O(N__20084),
            .I(rst));
    Odrv12 I__4601 (
            .O(N__20079),
            .I(rst));
    Odrv4 I__4600 (
            .O(N__20076),
            .I(rst));
    InMux I__4599 (
            .O(N__20061),
            .I(N__20058));
    LocalMux I__4598 (
            .O(N__20058),
            .I(\Lab_UT.scctrl.next_state_3_0 ));
    InMux I__4597 (
            .O(N__20055),
            .I(N__20049));
    InMux I__4596 (
            .O(N__20054),
            .I(N__20046));
    InMux I__4595 (
            .O(N__20053),
            .I(N__20040));
    InMux I__4594 (
            .O(N__20052),
            .I(N__20040));
    LocalMux I__4593 (
            .O(N__20049),
            .I(N__20034));
    LocalMux I__4592 (
            .O(N__20046),
            .I(N__20031));
    InMux I__4591 (
            .O(N__20045),
            .I(N__20028));
    LocalMux I__4590 (
            .O(N__20040),
            .I(N__20025));
    InMux I__4589 (
            .O(N__20039),
            .I(N__20018));
    InMux I__4588 (
            .O(N__20038),
            .I(N__20018));
    InMux I__4587 (
            .O(N__20037),
            .I(N__20018));
    Span4Mux_s3_h I__4586 (
            .O(N__20034),
            .I(N__20011));
    Span4Mux_v I__4585 (
            .O(N__20031),
            .I(N__20006));
    LocalMux I__4584 (
            .O(N__20028),
            .I(N__20006));
    Span4Mux_h I__4583 (
            .O(N__20025),
            .I(N__20001));
    LocalMux I__4582 (
            .O(N__20018),
            .I(N__20001));
    InMux I__4581 (
            .O(N__20017),
            .I(N__19998));
    InMux I__4580 (
            .O(N__20016),
            .I(N__19991));
    InMux I__4579 (
            .O(N__20015),
            .I(N__19991));
    InMux I__4578 (
            .O(N__20014),
            .I(N__19991));
    Odrv4 I__4577 (
            .O(N__20011),
            .I(\Lab_UT.scctrl.next_stateZ0Z_1 ));
    Odrv4 I__4576 (
            .O(N__20006),
            .I(\Lab_UT.scctrl.next_stateZ0Z_1 ));
    Odrv4 I__4575 (
            .O(N__20001),
            .I(\Lab_UT.scctrl.next_stateZ0Z_1 ));
    LocalMux I__4574 (
            .O(N__19998),
            .I(\Lab_UT.scctrl.next_stateZ0Z_1 ));
    LocalMux I__4573 (
            .O(N__19991),
            .I(\Lab_UT.scctrl.next_stateZ0Z_1 ));
    CascadeMux I__4572 (
            .O(N__19980),
            .I(\Lab_UT.scctrl.next_state_1_i_i_a2_1_0_1_cascade_ ));
    InMux I__4571 (
            .O(N__19977),
            .I(N__19973));
    InMux I__4570 (
            .O(N__19976),
            .I(N__19970));
    LocalMux I__4569 (
            .O(N__19973),
            .I(N__19967));
    LocalMux I__4568 (
            .O(N__19970),
            .I(N__19964));
    Span4Mux_v I__4567 (
            .O(N__19967),
            .I(N__19959));
    Span4Mux_v I__4566 (
            .O(N__19964),
            .I(N__19959));
    Odrv4 I__4565 (
            .O(N__19959),
            .I(\Lab_UT.scctrl.next_state_rst_0_6 ));
    InMux I__4564 (
            .O(N__19956),
            .I(N__19953));
    LocalMux I__4563 (
            .O(N__19953),
            .I(N__19950));
    Odrv12 I__4562 (
            .O(N__19950),
            .I(\Lab_UT.scctrl.N_398 ));
    InMux I__4561 (
            .O(N__19947),
            .I(N__19936));
    InMux I__4560 (
            .O(N__19946),
            .I(N__19936));
    CascadeMux I__4559 (
            .O(N__19945),
            .I(N__19931));
    CascadeMux I__4558 (
            .O(N__19944),
            .I(N__19927));
    CascadeMux I__4557 (
            .O(N__19943),
            .I(N__19923));
    CascadeMux I__4556 (
            .O(N__19942),
            .I(N__19920));
    CascadeMux I__4555 (
            .O(N__19941),
            .I(N__19917));
    LocalMux I__4554 (
            .O(N__19936),
            .I(N__19914));
    InMux I__4553 (
            .O(N__19935),
            .I(N__19911));
    CascadeMux I__4552 (
            .O(N__19934),
            .I(N__19908));
    InMux I__4551 (
            .O(N__19931),
            .I(N__19903));
    InMux I__4550 (
            .O(N__19930),
            .I(N__19900));
    InMux I__4549 (
            .O(N__19927),
            .I(N__19891));
    InMux I__4548 (
            .O(N__19926),
            .I(N__19891));
    InMux I__4547 (
            .O(N__19923),
            .I(N__19891));
    InMux I__4546 (
            .O(N__19920),
            .I(N__19891));
    InMux I__4545 (
            .O(N__19917),
            .I(N__19887));
    Span4Mux_v I__4544 (
            .O(N__19914),
            .I(N__19882));
    LocalMux I__4543 (
            .O(N__19911),
            .I(N__19882));
    InMux I__4542 (
            .O(N__19908),
            .I(N__19877));
    InMux I__4541 (
            .O(N__19907),
            .I(N__19877));
    CascadeMux I__4540 (
            .O(N__19906),
            .I(N__19874));
    LocalMux I__4539 (
            .O(N__19903),
            .I(N__19870));
    LocalMux I__4538 (
            .O(N__19900),
            .I(N__19865));
    LocalMux I__4537 (
            .O(N__19891),
            .I(N__19865));
    InMux I__4536 (
            .O(N__19890),
            .I(N__19862));
    LocalMux I__4535 (
            .O(N__19887),
            .I(N__19859));
    Span4Mux_v I__4534 (
            .O(N__19882),
            .I(N__19854));
    LocalMux I__4533 (
            .O(N__19877),
            .I(N__19854));
    InMux I__4532 (
            .O(N__19874),
            .I(N__19851));
    CascadeMux I__4531 (
            .O(N__19873),
            .I(N__19848));
    Span4Mux_v I__4530 (
            .O(N__19870),
            .I(N__19836));
    Span4Mux_h I__4529 (
            .O(N__19865),
            .I(N__19836));
    LocalMux I__4528 (
            .O(N__19862),
            .I(N__19836));
    Span4Mux_v I__4527 (
            .O(N__19859),
            .I(N__19836));
    Span4Mux_h I__4526 (
            .O(N__19854),
            .I(N__19836));
    LocalMux I__4525 (
            .O(N__19851),
            .I(N__19833));
    InMux I__4524 (
            .O(N__19848),
            .I(N__19828));
    InMux I__4523 (
            .O(N__19847),
            .I(N__19828));
    Span4Mux_v I__4522 (
            .O(N__19836),
            .I(N__19825));
    Span12Mux_s5_v I__4521 (
            .O(N__19833),
            .I(N__19822));
    LocalMux I__4520 (
            .O(N__19828),
            .I(\Lab_UT.scctrl.N_235_i_0 ));
    Odrv4 I__4519 (
            .O(N__19825),
            .I(\Lab_UT.scctrl.N_235_i_0 ));
    Odrv12 I__4518 (
            .O(N__19822),
            .I(\Lab_UT.scctrl.N_235_i_0 ));
    InMux I__4517 (
            .O(N__19815),
            .I(N__19810));
    InMux I__4516 (
            .O(N__19814),
            .I(N__19807));
    InMux I__4515 (
            .O(N__19813),
            .I(N__19804));
    LocalMux I__4514 (
            .O(N__19810),
            .I(N__19801));
    LocalMux I__4513 (
            .O(N__19807),
            .I(N__19796));
    LocalMux I__4512 (
            .O(N__19804),
            .I(N__19796));
    Span4Mux_s3_h I__4511 (
            .O(N__19801),
            .I(N__19793));
    Odrv12 I__4510 (
            .O(N__19796),
            .I(\Lab_UT.scctrl.N_240 ));
    Odrv4 I__4509 (
            .O(N__19793),
            .I(\Lab_UT.scctrl.N_240 ));
    CascadeMux I__4508 (
            .O(N__19788),
            .I(N__19785));
    InMux I__4507 (
            .O(N__19785),
            .I(N__19782));
    LocalMux I__4506 (
            .O(N__19782),
            .I(N__19779));
    Span4Mux_s2_h I__4505 (
            .O(N__19779),
            .I(N__19776));
    Span4Mux_v I__4504 (
            .O(N__19776),
            .I(N__19773));
    Odrv4 I__4503 (
            .O(N__19773),
            .I(\Lab_UT.scctrl.N_296 ));
    InMux I__4502 (
            .O(N__19770),
            .I(N__19767));
    LocalMux I__4501 (
            .O(N__19767),
            .I(N__19764));
    Odrv12 I__4500 (
            .O(N__19764),
            .I(\Lab_UT.scctrl.state_1_ret_1_RNICEVZ0Z81 ));
    CascadeMux I__4499 (
            .O(N__19761),
            .I(\Lab_UT.scctrl.G_24_i_1_cascade_ ));
    InMux I__4498 (
            .O(N__19758),
            .I(N__19755));
    LocalMux I__4497 (
            .O(N__19755),
            .I(N__19752));
    Odrv12 I__4496 (
            .O(N__19752),
            .I(\Lab_UT.scctrl.N_13_2 ));
    InMux I__4495 (
            .O(N__19749),
            .I(N__19745));
    InMux I__4494 (
            .O(N__19748),
            .I(N__19742));
    LocalMux I__4493 (
            .O(N__19745),
            .I(N__19737));
    LocalMux I__4492 (
            .O(N__19742),
            .I(N__19737));
    Span4Mux_h I__4491 (
            .O(N__19737),
            .I(N__19734));
    Odrv4 I__4490 (
            .O(N__19734),
            .I(\Lab_UT.scctrl.rst_retZ0 ));
    InMux I__4489 (
            .O(N__19731),
            .I(N__19722));
    CascadeMux I__4488 (
            .O(N__19730),
            .I(N__19719));
    InMux I__4487 (
            .O(N__19729),
            .I(N__19716));
    InMux I__4486 (
            .O(N__19728),
            .I(N__19713));
    InMux I__4485 (
            .O(N__19727),
            .I(N__19709));
    InMux I__4484 (
            .O(N__19726),
            .I(N__19706));
    InMux I__4483 (
            .O(N__19725),
            .I(N__19703));
    LocalMux I__4482 (
            .O(N__19722),
            .I(N__19700));
    InMux I__4481 (
            .O(N__19719),
            .I(N__19697));
    LocalMux I__4480 (
            .O(N__19716),
            .I(N__19694));
    LocalMux I__4479 (
            .O(N__19713),
            .I(N__19691));
    InMux I__4478 (
            .O(N__19712),
            .I(N__19688));
    LocalMux I__4477 (
            .O(N__19709),
            .I(N__19682));
    LocalMux I__4476 (
            .O(N__19706),
            .I(N__19682));
    LocalMux I__4475 (
            .O(N__19703),
            .I(N__19676));
    Span4Mux_v I__4474 (
            .O(N__19700),
            .I(N__19676));
    LocalMux I__4473 (
            .O(N__19697),
            .I(N__19671));
    Span4Mux_h I__4472 (
            .O(N__19694),
            .I(N__19671));
    Span4Mux_h I__4471 (
            .O(N__19691),
            .I(N__19664));
    LocalMux I__4470 (
            .O(N__19688),
            .I(N__19664));
    InMux I__4469 (
            .O(N__19687),
            .I(N__19661));
    Span4Mux_s2_h I__4468 (
            .O(N__19682),
            .I(N__19658));
    InMux I__4467 (
            .O(N__19681),
            .I(N__19655));
    Span4Mux_h I__4466 (
            .O(N__19676),
            .I(N__19650));
    Span4Mux_v I__4465 (
            .O(N__19671),
            .I(N__19650));
    InMux I__4464 (
            .O(N__19670),
            .I(N__19645));
    InMux I__4463 (
            .O(N__19669),
            .I(N__19645));
    Odrv4 I__4462 (
            .O(N__19664),
            .I(\Lab_UT.scctrl.state_i_2_2 ));
    LocalMux I__4461 (
            .O(N__19661),
            .I(\Lab_UT.scctrl.state_i_2_2 ));
    Odrv4 I__4460 (
            .O(N__19658),
            .I(\Lab_UT.scctrl.state_i_2_2 ));
    LocalMux I__4459 (
            .O(N__19655),
            .I(\Lab_UT.scctrl.state_i_2_2 ));
    Odrv4 I__4458 (
            .O(N__19650),
            .I(\Lab_UT.scctrl.state_i_2_2 ));
    LocalMux I__4457 (
            .O(N__19645),
            .I(\Lab_UT.scctrl.state_i_2_2 ));
    CascadeMux I__4456 (
            .O(N__19632),
            .I(\Lab_UT.scctrl.N_12_cascade_ ));
    InMux I__4455 (
            .O(N__19629),
            .I(N__19626));
    LocalMux I__4454 (
            .O(N__19626),
            .I(N__19623));
    Odrv12 I__4453 (
            .O(N__19623),
            .I(\Lab_UT.scctrl.N_8_0 ));
    InMux I__4452 (
            .O(N__19620),
            .I(N__19617));
    LocalMux I__4451 (
            .O(N__19617),
            .I(N__19614));
    Span4Mux_h I__4450 (
            .O(N__19614),
            .I(N__19611));
    Odrv4 I__4449 (
            .O(N__19611),
            .I(\Lab_UT.scctrl.g0_9_a2_4 ));
    CascadeMux I__4448 (
            .O(N__19608),
            .I(N__19604));
    InMux I__4447 (
            .O(N__19607),
            .I(N__19600));
    InMux I__4446 (
            .O(N__19604),
            .I(N__19591));
    InMux I__4445 (
            .O(N__19603),
            .I(N__19591));
    LocalMux I__4444 (
            .O(N__19600),
            .I(N__19588));
    InMux I__4443 (
            .O(N__19599),
            .I(N__19581));
    InMux I__4442 (
            .O(N__19598),
            .I(N__19581));
    InMux I__4441 (
            .O(N__19597),
            .I(N__19581));
    InMux I__4440 (
            .O(N__19596),
            .I(N__19578));
    LocalMux I__4439 (
            .O(N__19591),
            .I(N__19574));
    Span4Mux_v I__4438 (
            .O(N__19588),
            .I(N__19567));
    LocalMux I__4437 (
            .O(N__19581),
            .I(N__19567));
    LocalMux I__4436 (
            .O(N__19578),
            .I(N__19564));
    InMux I__4435 (
            .O(N__19577),
            .I(N__19561));
    Span4Mux_h I__4434 (
            .O(N__19574),
            .I(N__19558));
    InMux I__4433 (
            .O(N__19573),
            .I(N__19553));
    InMux I__4432 (
            .O(N__19572),
            .I(N__19553));
    Odrv4 I__4431 (
            .O(N__19567),
            .I(\Lab_UT.scctrl.state_3_rep1 ));
    Odrv4 I__4430 (
            .O(N__19564),
            .I(\Lab_UT.scctrl.state_3_rep1 ));
    LocalMux I__4429 (
            .O(N__19561),
            .I(\Lab_UT.scctrl.state_3_rep1 ));
    Odrv4 I__4428 (
            .O(N__19558),
            .I(\Lab_UT.scctrl.state_3_rep1 ));
    LocalMux I__4427 (
            .O(N__19553),
            .I(\Lab_UT.scctrl.state_3_rep1 ));
    InMux I__4426 (
            .O(N__19542),
            .I(N__19539));
    LocalMux I__4425 (
            .O(N__19539),
            .I(\Lab_UT.scctrl.g0_9_a3_0_0 ));
    CascadeMux I__4424 (
            .O(N__19536),
            .I(N__19531));
    CascadeMux I__4423 (
            .O(N__19535),
            .I(N__19526));
    CascadeMux I__4422 (
            .O(N__19534),
            .I(N__19522));
    InMux I__4421 (
            .O(N__19531),
            .I(N__19513));
    InMux I__4420 (
            .O(N__19530),
            .I(N__19513));
    InMux I__4419 (
            .O(N__19529),
            .I(N__19500));
    InMux I__4418 (
            .O(N__19526),
            .I(N__19500));
    InMux I__4417 (
            .O(N__19525),
            .I(N__19500));
    InMux I__4416 (
            .O(N__19522),
            .I(N__19500));
    InMux I__4415 (
            .O(N__19521),
            .I(N__19500));
    InMux I__4414 (
            .O(N__19520),
            .I(N__19500));
    InMux I__4413 (
            .O(N__19519),
            .I(N__19497));
    InMux I__4412 (
            .O(N__19518),
            .I(N__19489));
    LocalMux I__4411 (
            .O(N__19513),
            .I(N__19484));
    LocalMux I__4410 (
            .O(N__19500),
            .I(N__19484));
    LocalMux I__4409 (
            .O(N__19497),
            .I(N__19481));
    InMux I__4408 (
            .O(N__19496),
            .I(N__19476));
    InMux I__4407 (
            .O(N__19495),
            .I(N__19476));
    InMux I__4406 (
            .O(N__19494),
            .I(N__19473));
    InMux I__4405 (
            .O(N__19493),
            .I(N__19470));
    InMux I__4404 (
            .O(N__19492),
            .I(N__19467));
    LocalMux I__4403 (
            .O(N__19489),
            .I(N__19464));
    Span4Mux_v I__4402 (
            .O(N__19484),
            .I(N__19457));
    Span4Mux_s3_h I__4401 (
            .O(N__19481),
            .I(N__19457));
    LocalMux I__4400 (
            .O(N__19476),
            .I(N__19457));
    LocalMux I__4399 (
            .O(N__19473),
            .I(N__19454));
    LocalMux I__4398 (
            .O(N__19470),
            .I(N__19451));
    LocalMux I__4397 (
            .O(N__19467),
            .I(N__19444));
    Span4Mux_s3_h I__4396 (
            .O(N__19464),
            .I(N__19444));
    Span4Mux_v I__4395 (
            .O(N__19457),
            .I(N__19444));
    Span12Mux_s10_v I__4394 (
            .O(N__19454),
            .I(N__19441));
    Odrv12 I__4393 (
            .O(N__19451),
            .I(\Lab_UT.scctrl.next_stateZ0Z_3 ));
    Odrv4 I__4392 (
            .O(N__19444),
            .I(\Lab_UT.scctrl.next_stateZ0Z_3 ));
    Odrv12 I__4391 (
            .O(N__19441),
            .I(\Lab_UT.scctrl.next_stateZ0Z_3 ));
    InMux I__4390 (
            .O(N__19434),
            .I(N__19430));
    InMux I__4389 (
            .O(N__19433),
            .I(N__19427));
    LocalMux I__4388 (
            .O(N__19430),
            .I(N__19424));
    LocalMux I__4387 (
            .O(N__19427),
            .I(N__19421));
    Span4Mux_h I__4386 (
            .O(N__19424),
            .I(N__19418));
    Span4Mux_s2_h I__4385 (
            .O(N__19421),
            .I(N__19415));
    Odrv4 I__4384 (
            .O(N__19418),
            .I(\Lab_UT.scctrl.next_state_0_1 ));
    Odrv4 I__4383 (
            .O(N__19415),
            .I(\Lab_UT.scctrl.next_state_0_1 ));
    CascadeMux I__4382 (
            .O(N__19410),
            .I(\Lab_UT.scctrl.m90_i_o6_0_0_cascade_ ));
    InMux I__4381 (
            .O(N__19407),
            .I(N__19404));
    LocalMux I__4380 (
            .O(N__19404),
            .I(N__19401));
    Span4Mux_v I__4379 (
            .O(N__19401),
            .I(N__19398));
    Span4Mux_s1_h I__4378 (
            .O(N__19398),
            .I(N__19395));
    Odrv4 I__4377 (
            .O(N__19395),
            .I(\Lab_UT.scctrl.N_404_1 ));
    InMux I__4376 (
            .O(N__19392),
            .I(N__19386));
    InMux I__4375 (
            .O(N__19391),
            .I(N__19383));
    InMux I__4374 (
            .O(N__19390),
            .I(N__19380));
    InMux I__4373 (
            .O(N__19389),
            .I(N__19377));
    LocalMux I__4372 (
            .O(N__19386),
            .I(N__19373));
    LocalMux I__4371 (
            .O(N__19383),
            .I(N__19370));
    LocalMux I__4370 (
            .O(N__19380),
            .I(N__19366));
    LocalMux I__4369 (
            .O(N__19377),
            .I(N__19363));
    InMux I__4368 (
            .O(N__19376),
            .I(N__19360));
    Span4Mux_v I__4367 (
            .O(N__19373),
            .I(N__19355));
    Span4Mux_h I__4366 (
            .O(N__19370),
            .I(N__19355));
    InMux I__4365 (
            .O(N__19369),
            .I(N__19352));
    Odrv12 I__4364 (
            .O(N__19366),
            .I(\Lab_UT.scctrl.N_401 ));
    Odrv4 I__4363 (
            .O(N__19363),
            .I(\Lab_UT.scctrl.N_401 ));
    LocalMux I__4362 (
            .O(N__19360),
            .I(\Lab_UT.scctrl.N_401 ));
    Odrv4 I__4361 (
            .O(N__19355),
            .I(\Lab_UT.scctrl.N_401 ));
    LocalMux I__4360 (
            .O(N__19352),
            .I(\Lab_UT.scctrl.N_401 ));
    InMux I__4359 (
            .O(N__19341),
            .I(N__19337));
    InMux I__4358 (
            .O(N__19340),
            .I(N__19334));
    LocalMux I__4357 (
            .O(N__19337),
            .I(N__19328));
    LocalMux I__4356 (
            .O(N__19334),
            .I(N__19325));
    InMux I__4355 (
            .O(N__19333),
            .I(N__19322));
    InMux I__4354 (
            .O(N__19332),
            .I(N__19317));
    InMux I__4353 (
            .O(N__19331),
            .I(N__19317));
    Span4Mux_h I__4352 (
            .O(N__19328),
            .I(N__19312));
    Span4Mux_h I__4351 (
            .O(N__19325),
            .I(N__19309));
    LocalMux I__4350 (
            .O(N__19322),
            .I(N__19304));
    LocalMux I__4349 (
            .O(N__19317),
            .I(N__19304));
    InMux I__4348 (
            .O(N__19316),
            .I(N__19301));
    InMux I__4347 (
            .O(N__19315),
            .I(N__19298));
    Odrv4 I__4346 (
            .O(N__19312),
            .I(\Lab_UT.scctrl.N_399 ));
    Odrv4 I__4345 (
            .O(N__19309),
            .I(\Lab_UT.scctrl.N_399 ));
    Odrv12 I__4344 (
            .O(N__19304),
            .I(\Lab_UT.scctrl.N_399 ));
    LocalMux I__4343 (
            .O(N__19301),
            .I(\Lab_UT.scctrl.N_399 ));
    LocalMux I__4342 (
            .O(N__19298),
            .I(\Lab_UT.scctrl.N_399 ));
    CascadeMux I__4341 (
            .O(N__19287),
            .I(\Lab_UT.scctrl.g0_2_2_cascade_ ));
    InMux I__4340 (
            .O(N__19284),
            .I(N__19281));
    LocalMux I__4339 (
            .O(N__19281),
            .I(N__19278));
    Span4Mux_v I__4338 (
            .O(N__19278),
            .I(N__19275));
    Odrv4 I__4337 (
            .O(N__19275),
            .I(\Lab_UT.scctrl.g0_2_3 ));
    InMux I__4336 (
            .O(N__19272),
            .I(N__19269));
    LocalMux I__4335 (
            .O(N__19269),
            .I(N__19265));
    InMux I__4334 (
            .O(N__19268),
            .I(N__19262));
    Span4Mux_s2_h I__4333 (
            .O(N__19265),
            .I(N__19259));
    LocalMux I__4332 (
            .O(N__19262),
            .I(N__19256));
    Odrv4 I__4331 (
            .O(N__19259),
            .I(\Lab_UT.scctrl.g0_1_3 ));
    Odrv4 I__4330 (
            .O(N__19256),
            .I(\Lab_UT.scctrl.g0_1_3 ));
    InMux I__4329 (
            .O(N__19251),
            .I(N__19248));
    LocalMux I__4328 (
            .O(N__19248),
            .I(N__19238));
    InMux I__4327 (
            .O(N__19247),
            .I(N__19235));
    InMux I__4326 (
            .O(N__19246),
            .I(N__19222));
    InMux I__4325 (
            .O(N__19245),
            .I(N__19222));
    InMux I__4324 (
            .O(N__19244),
            .I(N__19222));
    InMux I__4323 (
            .O(N__19243),
            .I(N__19222));
    InMux I__4322 (
            .O(N__19242),
            .I(N__19222));
    InMux I__4321 (
            .O(N__19241),
            .I(N__19222));
    Odrv4 I__4320 (
            .O(N__19238),
            .I(\Lab_UT.scctrl.next_state_rst_2_2 ));
    LocalMux I__4319 (
            .O(N__19235),
            .I(\Lab_UT.scctrl.next_state_rst_2_2 ));
    LocalMux I__4318 (
            .O(N__19222),
            .I(\Lab_UT.scctrl.next_state_rst_2_2 ));
    InMux I__4317 (
            .O(N__19215),
            .I(N__19212));
    LocalMux I__4316 (
            .O(N__19212),
            .I(\Lab_UT.scctrl.N_13 ));
    InMux I__4315 (
            .O(N__19209),
            .I(N__19206));
    LocalMux I__4314 (
            .O(N__19206),
            .I(N__19203));
    Span4Mux_v I__4313 (
            .O(N__19203),
            .I(N__19200));
    Span4Mux_h I__4312 (
            .O(N__19200),
            .I(N__19197));
    Span4Mux_h I__4311 (
            .O(N__19197),
            .I(N__19194));
    Odrv4 I__4310 (
            .O(N__19194),
            .I(\Lab_UT.scctrl.N_404_0 ));
    CascadeMux I__4309 (
            .O(N__19191),
            .I(\Lab_UT.scctrl.N_5_3_cascade_ ));
    InMux I__4308 (
            .O(N__19188),
            .I(N__19185));
    LocalMux I__4307 (
            .O(N__19185),
            .I(N__19182));
    Odrv4 I__4306 (
            .O(N__19182),
            .I(\Lab_UT.scctrl.N_12_0 ));
    CascadeMux I__4305 (
            .O(N__19179),
            .I(N__19176));
    InMux I__4304 (
            .O(N__19176),
            .I(N__19173));
    LocalMux I__4303 (
            .O(N__19173),
            .I(N__19170));
    Span4Mux_s2_h I__4302 (
            .O(N__19170),
            .I(N__19167));
    Odrv4 I__4301 (
            .O(N__19167),
            .I(\Lab_UT.scctrl.G_18_i_a9_0 ));
    InMux I__4300 (
            .O(N__19164),
            .I(N__19161));
    LocalMux I__4299 (
            .O(N__19161),
            .I(\Lab_UT.scctrl.N_14_0 ));
    InMux I__4298 (
            .O(N__19158),
            .I(N__19148));
    CascadeMux I__4297 (
            .O(N__19157),
            .I(N__19145));
    CascadeMux I__4296 (
            .O(N__19156),
            .I(N__19141));
    InMux I__4295 (
            .O(N__19155),
            .I(N__19134));
    InMux I__4294 (
            .O(N__19154),
            .I(N__19134));
    InMux I__4293 (
            .O(N__19153),
            .I(N__19134));
    InMux I__4292 (
            .O(N__19152),
            .I(N__19126));
    InMux I__4291 (
            .O(N__19151),
            .I(N__19126));
    LocalMux I__4290 (
            .O(N__19148),
            .I(N__19122));
    InMux I__4289 (
            .O(N__19145),
            .I(N__19117));
    InMux I__4288 (
            .O(N__19144),
            .I(N__19117));
    InMux I__4287 (
            .O(N__19141),
            .I(N__19114));
    LocalMux I__4286 (
            .O(N__19134),
            .I(N__19111));
    InMux I__4285 (
            .O(N__19133),
            .I(N__19108));
    InMux I__4284 (
            .O(N__19132),
            .I(N__19105));
    InMux I__4283 (
            .O(N__19131),
            .I(N__19100));
    LocalMux I__4282 (
            .O(N__19126),
            .I(N__19097));
    InMux I__4281 (
            .O(N__19125),
            .I(N__19094));
    Span4Mux_v I__4280 (
            .O(N__19122),
            .I(N__19085));
    LocalMux I__4279 (
            .O(N__19117),
            .I(N__19085));
    LocalMux I__4278 (
            .O(N__19114),
            .I(N__19085));
    Span4Mux_v I__4277 (
            .O(N__19111),
            .I(N__19085));
    LocalMux I__4276 (
            .O(N__19108),
            .I(N__19082));
    LocalMux I__4275 (
            .O(N__19105),
            .I(N__19079));
    InMux I__4274 (
            .O(N__19104),
            .I(N__19074));
    InMux I__4273 (
            .O(N__19103),
            .I(N__19074));
    LocalMux I__4272 (
            .O(N__19100),
            .I(N__19071));
    Span4Mux_v I__4271 (
            .O(N__19097),
            .I(N__19068));
    LocalMux I__4270 (
            .O(N__19094),
            .I(N__19065));
    Span4Mux_v I__4269 (
            .O(N__19085),
            .I(N__19062));
    Span4Mux_v I__4268 (
            .O(N__19082),
            .I(N__19059));
    Sp12to4 I__4267 (
            .O(N__19079),
            .I(N__19054));
    LocalMux I__4266 (
            .O(N__19074),
            .I(N__19054));
    Span4Mux_s3_v I__4265 (
            .O(N__19071),
            .I(N__19049));
    Span4Mux_v I__4264 (
            .O(N__19068),
            .I(N__19049));
    Span4Mux_v I__4263 (
            .O(N__19065),
            .I(N__19042));
    Span4Mux_v I__4262 (
            .O(N__19062),
            .I(N__19042));
    Span4Mux_s0_h I__4261 (
            .O(N__19059),
            .I(N__19042));
    Odrv12 I__4260 (
            .O(N__19054),
            .I(\Lab_UT.scctrl.stateZ0Z_2 ));
    Odrv4 I__4259 (
            .O(N__19049),
            .I(\Lab_UT.scctrl.stateZ0Z_2 ));
    Odrv4 I__4258 (
            .O(N__19042),
            .I(\Lab_UT.scctrl.stateZ0Z_2 ));
    CascadeMux I__4257 (
            .O(N__19035),
            .I(N__19032));
    InMux I__4256 (
            .O(N__19032),
            .I(N__19028));
    CascadeMux I__4255 (
            .O(N__19031),
            .I(N__19025));
    LocalMux I__4254 (
            .O(N__19028),
            .I(N__19022));
    InMux I__4253 (
            .O(N__19025),
            .I(N__19019));
    Span4Mux_s2_h I__4252 (
            .O(N__19022),
            .I(N__19016));
    LocalMux I__4251 (
            .O(N__19019),
            .I(N__19013));
    Odrv4 I__4250 (
            .O(N__19016),
            .I(\Lab_UT.scctrl.N_5 ));
    Odrv4 I__4249 (
            .O(N__19013),
            .I(\Lab_UT.scctrl.N_5 ));
    CascadeMux I__4248 (
            .O(N__19008),
            .I(N__19005));
    InMux I__4247 (
            .O(N__19005),
            .I(N__19002));
    LocalMux I__4246 (
            .O(N__19002),
            .I(N__18999));
    Span4Mux_h I__4245 (
            .O(N__18999),
            .I(N__18996));
    Odrv4 I__4244 (
            .O(N__18996),
            .I(\Lab_UT.scctrl.N_21_0 ));
    CascadeMux I__4243 (
            .O(N__18993),
            .I(\Lab_UT.scctrl.G_10_i_o7_0_cascade_ ));
    InMux I__4242 (
            .O(N__18990),
            .I(N__18987));
    LocalMux I__4241 (
            .O(N__18987),
            .I(N__18984));
    Span4Mux_s3_h I__4240 (
            .O(N__18984),
            .I(N__18981));
    Odrv4 I__4239 (
            .O(N__18981),
            .I(\Lab_UT.scctrl.G_24_i_a7_4_2 ));
    InMux I__4238 (
            .O(N__18978),
            .I(N__18975));
    LocalMux I__4237 (
            .O(N__18975),
            .I(\Lab_UT.scctrl.G_18_i_a9_0_2 ));
    InMux I__4236 (
            .O(N__18972),
            .I(N__18969));
    LocalMux I__4235 (
            .O(N__18969),
            .I(N__18966));
    Span4Mux_v I__4234 (
            .O(N__18966),
            .I(N__18963));
    Odrv4 I__4233 (
            .O(N__18963),
            .I(\Lab_UT.scctrl.G_18_i_1 ));
    CascadeMux I__4232 (
            .O(N__18960),
            .I(\Lab_UT.scctrl.G_18_i_2_cascade_ ));
    CascadeMux I__4231 (
            .O(N__18957),
            .I(\Lab_UT.scctrl.G_18_i_4_cascade_ ));
    CascadeMux I__4230 (
            .O(N__18954),
            .I(N__18951));
    InMux I__4229 (
            .O(N__18951),
            .I(N__18948));
    LocalMux I__4228 (
            .O(N__18948),
            .I(N__18945));
    Span4Mux_h I__4227 (
            .O(N__18945),
            .I(N__18942));
    Span4Mux_v I__4226 (
            .O(N__18942),
            .I(N__18939));
    Odrv4 I__4225 (
            .O(N__18939),
            .I(\Lab_UT.scctrl.N_8_0_0 ));
    InMux I__4224 (
            .O(N__18936),
            .I(N__18933));
    LocalMux I__4223 (
            .O(N__18933),
            .I(N__18930));
    Span4Mux_s3_h I__4222 (
            .O(N__18930),
            .I(N__18927));
    Odrv4 I__4221 (
            .O(N__18927),
            .I(\Lab_UT.scctrl.g0_2_3_0 ));
    InMux I__4220 (
            .O(N__18924),
            .I(N__18921));
    LocalMux I__4219 (
            .O(N__18921),
            .I(N__18918));
    Span4Mux_h I__4218 (
            .O(N__18918),
            .I(N__18915));
    Span4Mux_v I__4217 (
            .O(N__18915),
            .I(N__18912));
    Odrv4 I__4216 (
            .O(N__18912),
            .I(\Lab_UT.scctrl.g0_2_2_0 ));
    CascadeMux I__4215 (
            .O(N__18909),
            .I(\Lab_UT.scctrl.next_state_2_0_cascade_ ));
    InMux I__4214 (
            .O(N__18906),
            .I(N__18900));
    InMux I__4213 (
            .O(N__18905),
            .I(N__18894));
    InMux I__4212 (
            .O(N__18904),
            .I(N__18891));
    CascadeMux I__4211 (
            .O(N__18903),
            .I(N__18888));
    LocalMux I__4210 (
            .O(N__18900),
            .I(N__18884));
    InMux I__4209 (
            .O(N__18899),
            .I(N__18879));
    InMux I__4208 (
            .O(N__18898),
            .I(N__18879));
    InMux I__4207 (
            .O(N__18897),
            .I(N__18876));
    LocalMux I__4206 (
            .O(N__18894),
            .I(N__18873));
    LocalMux I__4205 (
            .O(N__18891),
            .I(N__18870));
    InMux I__4204 (
            .O(N__18888),
            .I(N__18865));
    InMux I__4203 (
            .O(N__18887),
            .I(N__18865));
    Span4Mux_v I__4202 (
            .O(N__18884),
            .I(N__18862));
    LocalMux I__4201 (
            .O(N__18879),
            .I(N__18858));
    LocalMux I__4200 (
            .O(N__18876),
            .I(N__18849));
    Span4Mux_h I__4199 (
            .O(N__18873),
            .I(N__18849));
    Span4Mux_v I__4198 (
            .O(N__18870),
            .I(N__18849));
    LocalMux I__4197 (
            .O(N__18865),
            .I(N__18849));
    Span4Mux_v I__4196 (
            .O(N__18862),
            .I(N__18846));
    InMux I__4195 (
            .O(N__18861),
            .I(N__18843));
    Span4Mux_h I__4194 (
            .O(N__18858),
            .I(N__18838));
    Span4Mux_h I__4193 (
            .O(N__18849),
            .I(N__18838));
    Odrv4 I__4192 (
            .O(N__18846),
            .I(\Lab_UT.scctrl.N_260_i_0 ));
    LocalMux I__4191 (
            .O(N__18843),
            .I(\Lab_UT.scctrl.N_260_i_0 ));
    Odrv4 I__4190 (
            .O(N__18838),
            .I(\Lab_UT.scctrl.N_260_i_0 ));
    CascadeMux I__4189 (
            .O(N__18831),
            .I(N__18828));
    InMux I__4188 (
            .O(N__18828),
            .I(N__18825));
    LocalMux I__4187 (
            .O(N__18825),
            .I(N__18822));
    Span4Mux_v I__4186 (
            .O(N__18822),
            .I(N__18819));
    Span4Mux_h I__4185 (
            .O(N__18819),
            .I(N__18816));
    Odrv4 I__4184 (
            .O(N__18816),
            .I(\Lab_UT.scctrl.N_404_4 ));
    InMux I__4183 (
            .O(N__18813),
            .I(N__18809));
    InMux I__4182 (
            .O(N__18812),
            .I(N__18805));
    LocalMux I__4181 (
            .O(N__18809),
            .I(N__18800));
    InMux I__4180 (
            .O(N__18808),
            .I(N__18797));
    LocalMux I__4179 (
            .O(N__18805),
            .I(N__18794));
    InMux I__4178 (
            .O(N__18804),
            .I(N__18789));
    InMux I__4177 (
            .O(N__18803),
            .I(N__18789));
    Span4Mux_h I__4176 (
            .O(N__18800),
            .I(N__18776));
    LocalMux I__4175 (
            .O(N__18797),
            .I(N__18773));
    Span4Mux_s3_h I__4174 (
            .O(N__18794),
            .I(N__18770));
    LocalMux I__4173 (
            .O(N__18789),
            .I(N__18767));
    InMux I__4172 (
            .O(N__18788),
            .I(N__18764));
    InMux I__4171 (
            .O(N__18787),
            .I(N__18757));
    InMux I__4170 (
            .O(N__18786),
            .I(N__18757));
    InMux I__4169 (
            .O(N__18785),
            .I(N__18757));
    InMux I__4168 (
            .O(N__18784),
            .I(N__18748));
    InMux I__4167 (
            .O(N__18783),
            .I(N__18748));
    InMux I__4166 (
            .O(N__18782),
            .I(N__18748));
    InMux I__4165 (
            .O(N__18781),
            .I(N__18743));
    InMux I__4164 (
            .O(N__18780),
            .I(N__18743));
    InMux I__4163 (
            .O(N__18779),
            .I(N__18740));
    Span4Mux_v I__4162 (
            .O(N__18776),
            .I(N__18731));
    Span4Mux_h I__4161 (
            .O(N__18773),
            .I(N__18731));
    Span4Mux_h I__4160 (
            .O(N__18770),
            .I(N__18731));
    Span4Mux_h I__4159 (
            .O(N__18767),
            .I(N__18731));
    LocalMux I__4158 (
            .O(N__18764),
            .I(N__18728));
    LocalMux I__4157 (
            .O(N__18757),
            .I(N__18725));
    InMux I__4156 (
            .O(N__18756),
            .I(N__18722));
    InMux I__4155 (
            .O(N__18755),
            .I(N__18719));
    LocalMux I__4154 (
            .O(N__18748),
            .I(bu_rx_data_5));
    LocalMux I__4153 (
            .O(N__18743),
            .I(bu_rx_data_5));
    LocalMux I__4152 (
            .O(N__18740),
            .I(bu_rx_data_5));
    Odrv4 I__4151 (
            .O(N__18731),
            .I(bu_rx_data_5));
    Odrv4 I__4150 (
            .O(N__18728),
            .I(bu_rx_data_5));
    Odrv4 I__4149 (
            .O(N__18725),
            .I(bu_rx_data_5));
    LocalMux I__4148 (
            .O(N__18722),
            .I(bu_rx_data_5));
    LocalMux I__4147 (
            .O(N__18719),
            .I(bu_rx_data_5));
    InMux I__4146 (
            .O(N__18702),
            .I(N__18699));
    LocalMux I__4145 (
            .O(N__18699),
            .I(N__18696));
    Span4Mux_h I__4144 (
            .O(N__18696),
            .I(N__18693));
    Odrv4 I__4143 (
            .O(N__18693),
            .I(\Lab_UT.scctrl.g0_1_1_1 ));
    CascadeMux I__4142 (
            .O(N__18690),
            .I(N__18671));
    CascadeMux I__4141 (
            .O(N__18689),
            .I(N__18661));
    InMux I__4140 (
            .O(N__18688),
            .I(N__18655));
    InMux I__4139 (
            .O(N__18687),
            .I(N__18652));
    InMux I__4138 (
            .O(N__18686),
            .I(N__18647));
    InMux I__4137 (
            .O(N__18685),
            .I(N__18647));
    InMux I__4136 (
            .O(N__18684),
            .I(N__18642));
    InMux I__4135 (
            .O(N__18683),
            .I(N__18642));
    InMux I__4134 (
            .O(N__18682),
            .I(N__18633));
    InMux I__4133 (
            .O(N__18681),
            .I(N__18633));
    InMux I__4132 (
            .O(N__18680),
            .I(N__18633));
    InMux I__4131 (
            .O(N__18679),
            .I(N__18633));
    InMux I__4130 (
            .O(N__18678),
            .I(N__18624));
    InMux I__4129 (
            .O(N__18677),
            .I(N__18624));
    InMux I__4128 (
            .O(N__18676),
            .I(N__18624));
    InMux I__4127 (
            .O(N__18675),
            .I(N__18624));
    InMux I__4126 (
            .O(N__18674),
            .I(N__18606));
    InMux I__4125 (
            .O(N__18671),
            .I(N__18606));
    InMux I__4124 (
            .O(N__18670),
            .I(N__18606));
    InMux I__4123 (
            .O(N__18669),
            .I(N__18606));
    InMux I__4122 (
            .O(N__18668),
            .I(N__18606));
    InMux I__4121 (
            .O(N__18667),
            .I(N__18606));
    InMux I__4120 (
            .O(N__18666),
            .I(N__18606));
    InMux I__4119 (
            .O(N__18665),
            .I(N__18606));
    InMux I__4118 (
            .O(N__18664),
            .I(N__18595));
    InMux I__4117 (
            .O(N__18661),
            .I(N__18595));
    InMux I__4116 (
            .O(N__18660),
            .I(N__18595));
    InMux I__4115 (
            .O(N__18659),
            .I(N__18595));
    InMux I__4114 (
            .O(N__18658),
            .I(N__18595));
    LocalMux I__4113 (
            .O(N__18655),
            .I(N__18590));
    LocalMux I__4112 (
            .O(N__18652),
            .I(N__18590));
    LocalMux I__4111 (
            .O(N__18647),
            .I(N__18587));
    LocalMux I__4110 (
            .O(N__18642),
            .I(N__18580));
    LocalMux I__4109 (
            .O(N__18633),
            .I(N__18580));
    LocalMux I__4108 (
            .O(N__18624),
            .I(N__18580));
    CascadeMux I__4107 (
            .O(N__18623),
            .I(N__18577));
    LocalMux I__4106 (
            .O(N__18606),
            .I(N__18571));
    LocalMux I__4105 (
            .O(N__18595),
            .I(N__18566));
    Span4Mux_s2_v I__4104 (
            .O(N__18590),
            .I(N__18566));
    Span4Mux_v I__4103 (
            .O(N__18587),
            .I(N__18561));
    Span4Mux_v I__4102 (
            .O(N__18580),
            .I(N__18561));
    InMux I__4101 (
            .O(N__18577),
            .I(N__18558));
    InMux I__4100 (
            .O(N__18576),
            .I(N__18551));
    InMux I__4099 (
            .O(N__18575),
            .I(N__18551));
    InMux I__4098 (
            .O(N__18574),
            .I(N__18551));
    Span4Mux_v I__4097 (
            .O(N__18571),
            .I(N__18546));
    Span4Mux_v I__4096 (
            .O(N__18566),
            .I(N__18546));
    Span4Mux_h I__4095 (
            .O(N__18561),
            .I(N__18543));
    LocalMux I__4094 (
            .O(N__18558),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    LocalMux I__4093 (
            .O(N__18551),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    Odrv4 I__4092 (
            .O(N__18546),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    Odrv4 I__4091 (
            .O(N__18543),
            .I(\Lab_UT.scdp.binVal_ValidD ));
    InMux I__4090 (
            .O(N__18534),
            .I(N__18526));
    InMux I__4089 (
            .O(N__18533),
            .I(N__18526));
    InMux I__4088 (
            .O(N__18532),
            .I(N__18521));
    InMux I__4087 (
            .O(N__18531),
            .I(N__18521));
    LocalMux I__4086 (
            .O(N__18526),
            .I(N__18518));
    LocalMux I__4085 (
            .O(N__18521),
            .I(N__18512));
    Span4Mux_h I__4084 (
            .O(N__18518),
            .I(N__18509));
    InMux I__4083 (
            .O(N__18517),
            .I(N__18506));
    InMux I__4082 (
            .O(N__18516),
            .I(N__18501));
    InMux I__4081 (
            .O(N__18515),
            .I(N__18501));
    Span4Mux_h I__4080 (
            .O(N__18512),
            .I(N__18496));
    Span4Mux_h I__4079 (
            .O(N__18509),
            .I(N__18496));
    LocalMux I__4078 (
            .O(N__18506),
            .I(\Lab_UT.scdp.binValD_3 ));
    LocalMux I__4077 (
            .O(N__18501),
            .I(\Lab_UT.scdp.binValD_3 ));
    Odrv4 I__4076 (
            .O(N__18496),
            .I(\Lab_UT.scdp.binValD_3 ));
    InMux I__4075 (
            .O(N__18489),
            .I(N__18485));
    InMux I__4074 (
            .O(N__18488),
            .I(N__18479));
    LocalMux I__4073 (
            .O(N__18485),
            .I(N__18476));
    InMux I__4072 (
            .O(N__18484),
            .I(N__18473));
    InMux I__4071 (
            .O(N__18483),
            .I(N__18468));
    InMux I__4070 (
            .O(N__18482),
            .I(N__18468));
    LocalMux I__4069 (
            .O(N__18479),
            .I(\Lab_UT.state_1_RNI2IGHH_0_0 ));
    Odrv4 I__4068 (
            .O(N__18476),
            .I(\Lab_UT.state_1_RNI2IGHH_0_0 ));
    LocalMux I__4067 (
            .O(N__18473),
            .I(\Lab_UT.state_1_RNI2IGHH_0_0 ));
    LocalMux I__4066 (
            .O(N__18468),
            .I(\Lab_UT.state_1_RNI2IGHH_0_0 ));
    InMux I__4065 (
            .O(N__18459),
            .I(N__18455));
    CascadeMux I__4064 (
            .O(N__18458),
            .I(N__18452));
    LocalMux I__4063 (
            .O(N__18455),
            .I(N__18449));
    InMux I__4062 (
            .O(N__18452),
            .I(N__18446));
    Odrv12 I__4061 (
            .O(N__18449),
            .I(\Lab_UT.scdp.key2_7 ));
    LocalMux I__4060 (
            .O(N__18446),
            .I(\Lab_UT.scdp.key2_7 ));
    CascadeMux I__4059 (
            .O(N__18441),
            .I(N__18434));
    CascadeMux I__4058 (
            .O(N__18440),
            .I(N__18424));
    CascadeMux I__4057 (
            .O(N__18439),
            .I(N__18421));
    InMux I__4056 (
            .O(N__18438),
            .I(N__18417));
    InMux I__4055 (
            .O(N__18437),
            .I(N__18413));
    InMux I__4054 (
            .O(N__18434),
            .I(N__18410));
    CascadeMux I__4053 (
            .O(N__18433),
            .I(N__18407));
    InMux I__4052 (
            .O(N__18432),
            .I(N__18399));
    InMux I__4051 (
            .O(N__18431),
            .I(N__18399));
    InMux I__4050 (
            .O(N__18430),
            .I(N__18399));
    CascadeMux I__4049 (
            .O(N__18429),
            .I(N__18396));
    InMux I__4048 (
            .O(N__18428),
            .I(N__18392));
    InMux I__4047 (
            .O(N__18427),
            .I(N__18387));
    InMux I__4046 (
            .O(N__18424),
            .I(N__18387));
    InMux I__4045 (
            .O(N__18421),
            .I(N__18382));
    InMux I__4044 (
            .O(N__18420),
            .I(N__18382));
    LocalMux I__4043 (
            .O(N__18417),
            .I(N__18379));
    InMux I__4042 (
            .O(N__18416),
            .I(N__18376));
    LocalMux I__4041 (
            .O(N__18413),
            .I(N__18371));
    LocalMux I__4040 (
            .O(N__18410),
            .I(N__18371));
    InMux I__4039 (
            .O(N__18407),
            .I(N__18366));
    InMux I__4038 (
            .O(N__18406),
            .I(N__18366));
    LocalMux I__4037 (
            .O(N__18399),
            .I(N__18363));
    InMux I__4036 (
            .O(N__18396),
            .I(N__18360));
    CascadeMux I__4035 (
            .O(N__18395),
            .I(N__18357));
    LocalMux I__4034 (
            .O(N__18392),
            .I(N__18352));
    LocalMux I__4033 (
            .O(N__18387),
            .I(N__18347));
    LocalMux I__4032 (
            .O(N__18382),
            .I(N__18347));
    Span4Mux_s3_v I__4031 (
            .O(N__18379),
            .I(N__18338));
    LocalMux I__4030 (
            .O(N__18376),
            .I(N__18338));
    Span4Mux_h I__4029 (
            .O(N__18371),
            .I(N__18338));
    LocalMux I__4028 (
            .O(N__18366),
            .I(N__18338));
    Span4Mux_v I__4027 (
            .O(N__18363),
            .I(N__18333));
    LocalMux I__4026 (
            .O(N__18360),
            .I(N__18333));
    InMux I__4025 (
            .O(N__18357),
            .I(N__18330));
    InMux I__4024 (
            .O(N__18356),
            .I(N__18327));
    CascadeMux I__4023 (
            .O(N__18355),
            .I(N__18324));
    Span4Mux_v I__4022 (
            .O(N__18352),
            .I(N__18321));
    Span4Mux_v I__4021 (
            .O(N__18347),
            .I(N__18318));
    Span4Mux_v I__4020 (
            .O(N__18338),
            .I(N__18315));
    Span4Mux_v I__4019 (
            .O(N__18333),
            .I(N__18312));
    LocalMux I__4018 (
            .O(N__18330),
            .I(N__18307));
    LocalMux I__4017 (
            .O(N__18327),
            .I(N__18307));
    InMux I__4016 (
            .O(N__18324),
            .I(N__18304));
    Sp12to4 I__4015 (
            .O(N__18321),
            .I(N__18301));
    Span4Mux_v I__4014 (
            .O(N__18318),
            .I(N__18296));
    Span4Mux_s3_h I__4013 (
            .O(N__18315),
            .I(N__18296));
    Span4Mux_s2_h I__4012 (
            .O(N__18312),
            .I(N__18291));
    Span4Mux_v I__4011 (
            .O(N__18307),
            .I(N__18291));
    LocalMux I__4010 (
            .O(N__18304),
            .I(\Lab_UT.scctrl.state_i_1_0 ));
    Odrv12 I__4009 (
            .O(N__18301),
            .I(\Lab_UT.scctrl.state_i_1_0 ));
    Odrv4 I__4008 (
            .O(N__18296),
            .I(\Lab_UT.scctrl.state_i_1_0 ));
    Odrv4 I__4007 (
            .O(N__18291),
            .I(\Lab_UT.scctrl.state_i_1_0 ));
    InMux I__4006 (
            .O(N__18282),
            .I(N__18279));
    LocalMux I__4005 (
            .O(N__18279),
            .I(N__18272));
    InMux I__4004 (
            .O(N__18278),
            .I(N__18269));
    CascadeMux I__4003 (
            .O(N__18277),
            .I(N__18266));
    InMux I__4002 (
            .O(N__18276),
            .I(N__18260));
    InMux I__4001 (
            .O(N__18275),
            .I(N__18256));
    Span4Mux_h I__4000 (
            .O(N__18272),
            .I(N__18251));
    LocalMux I__3999 (
            .O(N__18269),
            .I(N__18251));
    InMux I__3998 (
            .O(N__18266),
            .I(N__18248));
    InMux I__3997 (
            .O(N__18265),
            .I(N__18242));
    InMux I__3996 (
            .O(N__18264),
            .I(N__18239));
    InMux I__3995 (
            .O(N__18263),
            .I(N__18235));
    LocalMux I__3994 (
            .O(N__18260),
            .I(N__18232));
    CascadeMux I__3993 (
            .O(N__18259),
            .I(N__18227));
    LocalMux I__3992 (
            .O(N__18256),
            .I(N__18222));
    Span4Mux_v I__3991 (
            .O(N__18251),
            .I(N__18217));
    LocalMux I__3990 (
            .O(N__18248),
            .I(N__18217));
    InMux I__3989 (
            .O(N__18247),
            .I(N__18212));
    InMux I__3988 (
            .O(N__18246),
            .I(N__18212));
    InMux I__3987 (
            .O(N__18245),
            .I(N__18209));
    LocalMux I__3986 (
            .O(N__18242),
            .I(N__18204));
    LocalMux I__3985 (
            .O(N__18239),
            .I(N__18204));
    InMux I__3984 (
            .O(N__18238),
            .I(N__18200));
    LocalMux I__3983 (
            .O(N__18235),
            .I(N__18197));
    Span4Mux_s2_h I__3982 (
            .O(N__18232),
            .I(N__18194));
    InMux I__3981 (
            .O(N__18231),
            .I(N__18191));
    InMux I__3980 (
            .O(N__18230),
            .I(N__18182));
    InMux I__3979 (
            .O(N__18227),
            .I(N__18182));
    InMux I__3978 (
            .O(N__18226),
            .I(N__18182));
    InMux I__3977 (
            .O(N__18225),
            .I(N__18182));
    Span4Mux_h I__3976 (
            .O(N__18222),
            .I(N__18177));
    Span4Mux_h I__3975 (
            .O(N__18217),
            .I(N__18177));
    LocalMux I__3974 (
            .O(N__18212),
            .I(N__18174));
    LocalMux I__3973 (
            .O(N__18209),
            .I(N__18169));
    Span12Mux_v I__3972 (
            .O(N__18204),
            .I(N__18169));
    InMux I__3971 (
            .O(N__18203),
            .I(N__18166));
    LocalMux I__3970 (
            .O(N__18200),
            .I(\Lab_UT.scctrl.N_296_i_0 ));
    Odrv4 I__3969 (
            .O(N__18197),
            .I(\Lab_UT.scctrl.N_296_i_0 ));
    Odrv4 I__3968 (
            .O(N__18194),
            .I(\Lab_UT.scctrl.N_296_i_0 ));
    LocalMux I__3967 (
            .O(N__18191),
            .I(\Lab_UT.scctrl.N_296_i_0 ));
    LocalMux I__3966 (
            .O(N__18182),
            .I(\Lab_UT.scctrl.N_296_i_0 ));
    Odrv4 I__3965 (
            .O(N__18177),
            .I(\Lab_UT.scctrl.N_296_i_0 ));
    Odrv12 I__3964 (
            .O(N__18174),
            .I(\Lab_UT.scctrl.N_296_i_0 ));
    Odrv12 I__3963 (
            .O(N__18169),
            .I(\Lab_UT.scctrl.N_296_i_0 ));
    LocalMux I__3962 (
            .O(N__18166),
            .I(\Lab_UT.scctrl.N_296_i_0 ));
    InMux I__3961 (
            .O(N__18147),
            .I(N__18144));
    LocalMux I__3960 (
            .O(N__18144),
            .I(N__18141));
    Span4Mux_v I__3959 (
            .O(N__18141),
            .I(N__18138));
    Span4Mux_h I__3958 (
            .O(N__18138),
            .I(N__18135));
    Odrv4 I__3957 (
            .O(N__18135),
            .I(\Lab_UT.scctrl.next_state_RNO_1Z0Z_1 ));
    CascadeMux I__3956 (
            .O(N__18132),
            .I(\Lab_UT.scctrl.N_319_cascade_ ));
    InMux I__3955 (
            .O(N__18129),
            .I(N__18126));
    LocalMux I__3954 (
            .O(N__18126),
            .I(N__18123));
    Span4Mux_v I__3953 (
            .O(N__18123),
            .I(N__18120));
    Odrv4 I__3952 (
            .O(N__18120),
            .I(\Lab_UT.scctrl.next_state_rst_1_0 ));
    CascadeMux I__3951 (
            .O(N__18117),
            .I(\Lab_UT.scctrl.N_414_cascade_ ));
    InMux I__3950 (
            .O(N__18114),
            .I(N__18108));
    InMux I__3949 (
            .O(N__18113),
            .I(N__18108));
    LocalMux I__3948 (
            .O(N__18108),
            .I(N__18105));
    Span4Mux_v I__3947 (
            .O(N__18105),
            .I(N__18102));
    Odrv4 I__3946 (
            .O(N__18102),
            .I(\Lab_UT.scctrl.next_state_rst_1_2 ));
    InMux I__3945 (
            .O(N__18099),
            .I(N__18096));
    LocalMux I__3944 (
            .O(N__18096),
            .I(N__18093));
    Span4Mux_h I__3943 (
            .O(N__18093),
            .I(N__18090));
    Odrv4 I__3942 (
            .O(N__18090),
            .I(\Lab_UT.scctrl.N_319_1 ));
    CascadeMux I__3941 (
            .O(N__18087),
            .I(N__18082));
    CascadeMux I__3940 (
            .O(N__18086),
            .I(N__18079));
    CascadeMux I__3939 (
            .O(N__18085),
            .I(N__18076));
    InMux I__3938 (
            .O(N__18082),
            .I(N__18073));
    InMux I__3937 (
            .O(N__18079),
            .I(N__18068));
    InMux I__3936 (
            .O(N__18076),
            .I(N__18062));
    LocalMux I__3935 (
            .O(N__18073),
            .I(N__18059));
    InMux I__3934 (
            .O(N__18072),
            .I(N__18055));
    CascadeMux I__3933 (
            .O(N__18071),
            .I(N__18051));
    LocalMux I__3932 (
            .O(N__18068),
            .I(N__18048));
    InMux I__3931 (
            .O(N__18067),
            .I(N__18043));
    InMux I__3930 (
            .O(N__18066),
            .I(N__18043));
    InMux I__3929 (
            .O(N__18065),
            .I(N__18040));
    LocalMux I__3928 (
            .O(N__18062),
            .I(N__18035));
    Span4Mux_v I__3927 (
            .O(N__18059),
            .I(N__18032));
    CascadeMux I__3926 (
            .O(N__18058),
            .I(N__18029));
    LocalMux I__3925 (
            .O(N__18055),
            .I(N__18025));
    CascadeMux I__3924 (
            .O(N__18054),
            .I(N__18022));
    InMux I__3923 (
            .O(N__18051),
            .I(N__18019));
    Span4Mux_h I__3922 (
            .O(N__18048),
            .I(N__18014));
    LocalMux I__3921 (
            .O(N__18043),
            .I(N__18014));
    LocalMux I__3920 (
            .O(N__18040),
            .I(N__18011));
    InMux I__3919 (
            .O(N__18039),
            .I(N__18008));
    InMux I__3918 (
            .O(N__18038),
            .I(N__18005));
    Span4Mux_v I__3917 (
            .O(N__18035),
            .I(N__17999));
    Span4Mux_s3_h I__3916 (
            .O(N__18032),
            .I(N__17999));
    InMux I__3915 (
            .O(N__18029),
            .I(N__17994));
    InMux I__3914 (
            .O(N__18028),
            .I(N__17994));
    Span4Mux_s2_h I__3913 (
            .O(N__18025),
            .I(N__17991));
    InMux I__3912 (
            .O(N__18022),
            .I(N__17988));
    LocalMux I__3911 (
            .O(N__18019),
            .I(N__17983));
    Span4Mux_s3_h I__3910 (
            .O(N__18014),
            .I(N__17983));
    Span4Mux_v I__3909 (
            .O(N__18011),
            .I(N__17976));
    LocalMux I__3908 (
            .O(N__18008),
            .I(N__17976));
    LocalMux I__3907 (
            .O(N__18005),
            .I(N__17976));
    InMux I__3906 (
            .O(N__18004),
            .I(N__17973));
    Span4Mux_v I__3905 (
            .O(N__17999),
            .I(N__17968));
    LocalMux I__3904 (
            .O(N__17994),
            .I(N__17968));
    Odrv4 I__3903 (
            .O(N__17991),
            .I(\Lab_UT.scctrl.state_2_rep2 ));
    LocalMux I__3902 (
            .O(N__17988),
            .I(\Lab_UT.scctrl.state_2_rep2 ));
    Odrv4 I__3901 (
            .O(N__17983),
            .I(\Lab_UT.scctrl.state_2_rep2 ));
    Odrv4 I__3900 (
            .O(N__17976),
            .I(\Lab_UT.scctrl.state_2_rep2 ));
    LocalMux I__3899 (
            .O(N__17973),
            .I(\Lab_UT.scctrl.state_2_rep2 ));
    Odrv4 I__3898 (
            .O(N__17968),
            .I(\Lab_UT.scctrl.state_2_rep2 ));
    CascadeMux I__3897 (
            .O(N__17955),
            .I(\Lab_UT.scctrl.N_7_1_cascade_ ));
    InMux I__3896 (
            .O(N__17952),
            .I(N__17945));
    InMux I__3895 (
            .O(N__17951),
            .I(N__17936));
    InMux I__3894 (
            .O(N__17950),
            .I(N__17936));
    InMux I__3893 (
            .O(N__17949),
            .I(N__17936));
    InMux I__3892 (
            .O(N__17948),
            .I(N__17936));
    LocalMux I__3891 (
            .O(N__17945),
            .I(\Lab_UT.state_ret_12_RNIUVHQG_0 ));
    LocalMux I__3890 (
            .O(N__17936),
            .I(\Lab_UT.state_ret_12_RNIUVHQG_0 ));
    InMux I__3889 (
            .O(N__17931),
            .I(N__17927));
    CascadeMux I__3888 (
            .O(N__17930),
            .I(N__17924));
    LocalMux I__3887 (
            .O(N__17927),
            .I(N__17921));
    InMux I__3886 (
            .O(N__17924),
            .I(N__17918));
    Odrv12 I__3885 (
            .O(N__17921),
            .I(\Lab_UT.scdp.key3_3 ));
    LocalMux I__3884 (
            .O(N__17918),
            .I(\Lab_UT.scdp.key3_3 ));
    CascadeMux I__3883 (
            .O(N__17913),
            .I(N__17910));
    InMux I__3882 (
            .O(N__17910),
            .I(N__17906));
    InMux I__3881 (
            .O(N__17909),
            .I(N__17903));
    LocalMux I__3880 (
            .O(N__17906),
            .I(\Lab_UT.scdp.val_0_tz_3 ));
    LocalMux I__3879 (
            .O(N__17903),
            .I(\Lab_UT.scdp.val_0_tz_3 ));
    CascadeMux I__3878 (
            .O(N__17898),
            .I(N__17887));
    CascadeMux I__3877 (
            .O(N__17897),
            .I(N__17881));
    CascadeMux I__3876 (
            .O(N__17896),
            .I(N__17878));
    CascadeMux I__3875 (
            .O(N__17895),
            .I(N__17875));
    CascadeMux I__3874 (
            .O(N__17894),
            .I(N__17872));
    InMux I__3873 (
            .O(N__17893),
            .I(N__17869));
    InMux I__3872 (
            .O(N__17892),
            .I(N__17866));
    InMux I__3871 (
            .O(N__17891),
            .I(N__17859));
    InMux I__3870 (
            .O(N__17890),
            .I(N__17859));
    InMux I__3869 (
            .O(N__17887),
            .I(N__17859));
    InMux I__3868 (
            .O(N__17886),
            .I(N__17856));
    InMux I__3867 (
            .O(N__17885),
            .I(N__17852));
    InMux I__3866 (
            .O(N__17884),
            .I(N__17841));
    InMux I__3865 (
            .O(N__17881),
            .I(N__17841));
    InMux I__3864 (
            .O(N__17878),
            .I(N__17841));
    InMux I__3863 (
            .O(N__17875),
            .I(N__17841));
    InMux I__3862 (
            .O(N__17872),
            .I(N__17841));
    LocalMux I__3861 (
            .O(N__17869),
            .I(N__17834));
    LocalMux I__3860 (
            .O(N__17866),
            .I(N__17834));
    LocalMux I__3859 (
            .O(N__17859),
            .I(N__17834));
    LocalMux I__3858 (
            .O(N__17856),
            .I(N__17831));
    InMux I__3857 (
            .O(N__17855),
            .I(N__17828));
    LocalMux I__3856 (
            .O(N__17852),
            .I(N__17820));
    LocalMux I__3855 (
            .O(N__17841),
            .I(N__17820));
    Span4Mux_h I__3854 (
            .O(N__17834),
            .I(N__17820));
    Span4Mux_h I__3853 (
            .O(N__17831),
            .I(N__17817));
    LocalMux I__3852 (
            .O(N__17828),
            .I(N__17814));
    InMux I__3851 (
            .O(N__17827),
            .I(N__17811));
    Span4Mux_v I__3850 (
            .O(N__17820),
            .I(N__17808));
    Span4Mux_v I__3849 (
            .O(N__17817),
            .I(N__17801));
    Span4Mux_h I__3848 (
            .O(N__17814),
            .I(N__17801));
    LocalMux I__3847 (
            .O(N__17811),
            .I(N__17801));
    Span4Mux_h I__3846 (
            .O(N__17808),
            .I(N__17798));
    Odrv4 I__3845 (
            .O(N__17801),
            .I(bu_rx_data_i_2_3));
    Odrv4 I__3844 (
            .O(N__17798),
            .I(bu_rx_data_i_2_3));
    InMux I__3843 (
            .O(N__17793),
            .I(N__17788));
    InMux I__3842 (
            .O(N__17792),
            .I(N__17785));
    CascadeMux I__3841 (
            .O(N__17791),
            .I(N__17782));
    LocalMux I__3840 (
            .O(N__17788),
            .I(N__17779));
    LocalMux I__3839 (
            .O(N__17785),
            .I(N__17776));
    InMux I__3838 (
            .O(N__17782),
            .I(N__17773));
    Span4Mux_h I__3837 (
            .O(N__17779),
            .I(N__17768));
    Span4Mux_v I__3836 (
            .O(N__17776),
            .I(N__17768));
    LocalMux I__3835 (
            .O(N__17773),
            .I(\buart.Z_rx.N_301 ));
    Odrv4 I__3834 (
            .O(N__17768),
            .I(\buart.Z_rx.N_301 ));
    InMux I__3833 (
            .O(N__17763),
            .I(N__17759));
    InMux I__3832 (
            .O(N__17762),
            .I(N__17756));
    LocalMux I__3831 (
            .O(N__17759),
            .I(N__17753));
    LocalMux I__3830 (
            .O(N__17756),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    Odrv12 I__3829 (
            .O(N__17753),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    CascadeMux I__3828 (
            .O(N__17748),
            .I(N__17744));
    InMux I__3827 (
            .O(N__17747),
            .I(N__17736));
    InMux I__3826 (
            .O(N__17744),
            .I(N__17736));
    InMux I__3825 (
            .O(N__17743),
            .I(N__17736));
    LocalMux I__3824 (
            .O(N__17736),
            .I(N__17731));
    InMux I__3823 (
            .O(N__17735),
            .I(N__17728));
    InMux I__3822 (
            .O(N__17734),
            .I(N__17725));
    Span4Mux_v I__3821 (
            .O(N__17731),
            .I(N__17720));
    LocalMux I__3820 (
            .O(N__17728),
            .I(N__17720));
    LocalMux I__3819 (
            .O(N__17725),
            .I(N__17717));
    Span4Mux_h I__3818 (
            .O(N__17720),
            .I(N__17714));
    Span4Mux_h I__3817 (
            .O(N__17717),
            .I(N__17711));
    Span4Mux_v I__3816 (
            .O(N__17714),
            .I(N__17708));
    Odrv4 I__3815 (
            .O(N__17711),
            .I(buart__rx_hh_1));
    Odrv4 I__3814 (
            .O(N__17708),
            .I(buart__rx_hh_1));
    InMux I__3813 (
            .O(N__17703),
            .I(N__17691));
    InMux I__3812 (
            .O(N__17702),
            .I(N__17686));
    InMux I__3811 (
            .O(N__17701),
            .I(N__17686));
    CascadeMux I__3810 (
            .O(N__17700),
            .I(N__17682));
    CascadeMux I__3809 (
            .O(N__17699),
            .I(N__17679));
    CascadeMux I__3808 (
            .O(N__17698),
            .I(N__17676));
    InMux I__3807 (
            .O(N__17697),
            .I(N__17666));
    InMux I__3806 (
            .O(N__17696),
            .I(N__17666));
    InMux I__3805 (
            .O(N__17695),
            .I(N__17666));
    InMux I__3804 (
            .O(N__17694),
            .I(N__17666));
    LocalMux I__3803 (
            .O(N__17691),
            .I(N__17661));
    LocalMux I__3802 (
            .O(N__17686),
            .I(N__17661));
    InMux I__3801 (
            .O(N__17685),
            .I(N__17652));
    InMux I__3800 (
            .O(N__17682),
            .I(N__17652));
    InMux I__3799 (
            .O(N__17679),
            .I(N__17652));
    InMux I__3798 (
            .O(N__17676),
            .I(N__17652));
    InMux I__3797 (
            .O(N__17675),
            .I(N__17649));
    LocalMux I__3796 (
            .O(N__17666),
            .I(N__17646));
    Span4Mux_v I__3795 (
            .O(N__17661),
            .I(N__17641));
    LocalMux I__3794 (
            .O(N__17652),
            .I(N__17641));
    LocalMux I__3793 (
            .O(N__17649),
            .I(N__17634));
    Span4Mux_v I__3792 (
            .O(N__17646),
            .I(N__17634));
    Span4Mux_h I__3791 (
            .O(N__17641),
            .I(N__17634));
    Span4Mux_h I__3790 (
            .O(N__17634),
            .I(N__17631));
    Odrv4 I__3789 (
            .O(N__17631),
            .I(\buart.Z_rx.startbit ));
    InMux I__3788 (
            .O(N__17628),
            .I(N__17623));
    InMux I__3787 (
            .O(N__17627),
            .I(N__17618));
    InMux I__3786 (
            .O(N__17626),
            .I(N__17618));
    LocalMux I__3785 (
            .O(N__17623),
            .I(N__17610));
    LocalMux I__3784 (
            .O(N__17618),
            .I(N__17610));
    InMux I__3783 (
            .O(N__17617),
            .I(N__17605));
    InMux I__3782 (
            .O(N__17616),
            .I(N__17605));
    InMux I__3781 (
            .O(N__17615),
            .I(N__17602));
    Span4Mux_v I__3780 (
            .O(N__17610),
            .I(N__17597));
    LocalMux I__3779 (
            .O(N__17605),
            .I(N__17594));
    LocalMux I__3778 (
            .O(N__17602),
            .I(N__17591));
    InMux I__3777 (
            .O(N__17601),
            .I(N__17586));
    InMux I__3776 (
            .O(N__17600),
            .I(N__17586));
    Odrv4 I__3775 (
            .O(N__17597),
            .I(\Lab_UT.scdp.binValD_0 ));
    Odrv4 I__3774 (
            .O(N__17594),
            .I(\Lab_UT.scdp.binValD_0 ));
    Odrv4 I__3773 (
            .O(N__17591),
            .I(\Lab_UT.scdp.binValD_0 ));
    LocalMux I__3772 (
            .O(N__17586),
            .I(\Lab_UT.scdp.binValD_0 ));
    InMux I__3771 (
            .O(N__17577),
            .I(N__17574));
    LocalMux I__3770 (
            .O(N__17574),
            .I(N__17570));
    CascadeMux I__3769 (
            .O(N__17573),
            .I(N__17567));
    Span4Mux_v I__3768 (
            .O(N__17570),
            .I(N__17564));
    InMux I__3767 (
            .O(N__17567),
            .I(N__17561));
    Odrv4 I__3766 (
            .O(N__17564),
            .I(\Lab_UT.scdp.key0_0 ));
    LocalMux I__3765 (
            .O(N__17561),
            .I(\Lab_UT.scdp.key0_0 ));
    InMux I__3764 (
            .O(N__17556),
            .I(N__17550));
    InMux I__3763 (
            .O(N__17555),
            .I(N__17550));
    LocalMux I__3762 (
            .O(N__17550),
            .I(N__17546));
    InMux I__3761 (
            .O(N__17549),
            .I(N__17541));
    Span4Mux_h I__3760 (
            .O(N__17546),
            .I(N__17538));
    InMux I__3759 (
            .O(N__17545),
            .I(N__17533));
    InMux I__3758 (
            .O(N__17544),
            .I(N__17533));
    LocalMux I__3757 (
            .O(N__17541),
            .I(\Lab_UT.state_1_RNIO1RJH_0_2 ));
    Odrv4 I__3756 (
            .O(N__17538),
            .I(\Lab_UT.state_1_RNIO1RJH_0_2 ));
    LocalMux I__3755 (
            .O(N__17533),
            .I(\Lab_UT.state_1_RNIO1RJH_0_2 ));
    InMux I__3754 (
            .O(N__17526),
            .I(N__17522));
    CascadeMux I__3753 (
            .O(N__17525),
            .I(N__17519));
    LocalMux I__3752 (
            .O(N__17522),
            .I(N__17516));
    InMux I__3751 (
            .O(N__17519),
            .I(N__17513));
    Odrv12 I__3750 (
            .O(N__17516),
            .I(\Lab_UT.scdp.key0_1 ));
    LocalMux I__3749 (
            .O(N__17513),
            .I(\Lab_UT.scdp.key0_1 ));
    InMux I__3748 (
            .O(N__17508),
            .I(N__17501));
    InMux I__3747 (
            .O(N__17507),
            .I(N__17498));
    InMux I__3746 (
            .O(N__17506),
            .I(N__17493));
    InMux I__3745 (
            .O(N__17505),
            .I(N__17493));
    InMux I__3744 (
            .O(N__17504),
            .I(N__17490));
    LocalMux I__3743 (
            .O(N__17501),
            .I(\Lab_UT.state_1_ret_3_RNI23U7H_0 ));
    LocalMux I__3742 (
            .O(N__17498),
            .I(\Lab_UT.state_1_ret_3_RNI23U7H_0 ));
    LocalMux I__3741 (
            .O(N__17493),
            .I(\Lab_UT.state_1_ret_3_RNI23U7H_0 ));
    LocalMux I__3740 (
            .O(N__17490),
            .I(\Lab_UT.state_1_ret_3_RNI23U7H_0 ));
    InMux I__3739 (
            .O(N__17481),
            .I(N__17478));
    LocalMux I__3738 (
            .O(N__17478),
            .I(N__17475));
    Span4Mux_v I__3737 (
            .O(N__17475),
            .I(N__17471));
    CascadeMux I__3736 (
            .O(N__17474),
            .I(N__17468));
    Span4Mux_h I__3735 (
            .O(N__17471),
            .I(N__17465));
    InMux I__3734 (
            .O(N__17468),
            .I(N__17462));
    Odrv4 I__3733 (
            .O(N__17465),
            .I(\Lab_UT.scdp.key1_5 ));
    LocalMux I__3732 (
            .O(N__17462),
            .I(\Lab_UT.scdp.key1_5 ));
    InMux I__3731 (
            .O(N__17457),
            .I(N__17450));
    InMux I__3730 (
            .O(N__17456),
            .I(N__17447));
    InMux I__3729 (
            .O(N__17455),
            .I(N__17444));
    InMux I__3728 (
            .O(N__17454),
            .I(N__17439));
    InMux I__3727 (
            .O(N__17453),
            .I(N__17439));
    LocalMux I__3726 (
            .O(N__17450),
            .I(\Lab_UT.state_ret_RNIK5UKH_0 ));
    LocalMux I__3725 (
            .O(N__17447),
            .I(\Lab_UT.state_ret_RNIK5UKH_0 ));
    LocalMux I__3724 (
            .O(N__17444),
            .I(\Lab_UT.state_ret_RNIK5UKH_0 ));
    LocalMux I__3723 (
            .O(N__17439),
            .I(\Lab_UT.state_ret_RNIK5UKH_0 ));
    InMux I__3722 (
            .O(N__17430),
            .I(N__17427));
    LocalMux I__3721 (
            .O(N__17427),
            .I(N__17423));
    CascadeMux I__3720 (
            .O(N__17426),
            .I(N__17420));
    Span4Mux_h I__3719 (
            .O(N__17423),
            .I(N__17417));
    InMux I__3718 (
            .O(N__17420),
            .I(N__17414));
    Odrv4 I__3717 (
            .O(N__17417),
            .I(\Lab_UT.scdp.key2_3 ));
    LocalMux I__3716 (
            .O(N__17414),
            .I(\Lab_UT.scdp.key2_3 ));
    InMux I__3715 (
            .O(N__17409),
            .I(N__17403));
    InMux I__3714 (
            .O(N__17408),
            .I(N__17403));
    LocalMux I__3713 (
            .O(N__17403),
            .I(N__17399));
    InMux I__3712 (
            .O(N__17402),
            .I(N__17396));
    Span4Mux_v I__3711 (
            .O(N__17399),
            .I(N__17388));
    LocalMux I__3710 (
            .O(N__17396),
            .I(N__17388));
    InMux I__3709 (
            .O(N__17395),
            .I(N__17381));
    InMux I__3708 (
            .O(N__17394),
            .I(N__17381));
    InMux I__3707 (
            .O(N__17393),
            .I(N__17381));
    Span4Mux_h I__3706 (
            .O(N__17388),
            .I(N__17376));
    LocalMux I__3705 (
            .O(N__17381),
            .I(N__17376));
    Span4Mux_v I__3704 (
            .O(N__17376),
            .I(N__17371));
    InMux I__3703 (
            .O(N__17375),
            .I(N__17366));
    InMux I__3702 (
            .O(N__17374),
            .I(N__17366));
    Span4Mux_s3_h I__3701 (
            .O(N__17371),
            .I(N__17363));
    LocalMux I__3700 (
            .O(N__17366),
            .I(\Lab_UT.scdp.binValD_1 ));
    Odrv4 I__3699 (
            .O(N__17363),
            .I(\Lab_UT.scdp.binValD_1 ));
    InMux I__3698 (
            .O(N__17358),
            .I(N__17351));
    InMux I__3697 (
            .O(N__17357),
            .I(N__17348));
    InMux I__3696 (
            .O(N__17356),
            .I(N__17341));
    InMux I__3695 (
            .O(N__17355),
            .I(N__17341));
    InMux I__3694 (
            .O(N__17354),
            .I(N__17341));
    LocalMux I__3693 (
            .O(N__17351),
            .I(\Lab_UT.state_ret_12_RNI2SEPG_0 ));
    LocalMux I__3692 (
            .O(N__17348),
            .I(\Lab_UT.state_ret_12_RNI2SEPG_0 ));
    LocalMux I__3691 (
            .O(N__17341),
            .I(\Lab_UT.state_ret_12_RNI2SEPG_0 ));
    InMux I__3690 (
            .O(N__17334),
            .I(N__17331));
    LocalMux I__3689 (
            .O(N__17331),
            .I(N__17327));
    CascadeMux I__3688 (
            .O(N__17330),
            .I(N__17324));
    Span4Mux_s2_v I__3687 (
            .O(N__17327),
            .I(N__17321));
    InMux I__3686 (
            .O(N__17324),
            .I(N__17318));
    Odrv4 I__3685 (
            .O(N__17321),
            .I(\Lab_UT.scdp.key1_1 ));
    LocalMux I__3684 (
            .O(N__17318),
            .I(\Lab_UT.scdp.key1_1 ));
    CascadeMux I__3683 (
            .O(N__17313),
            .I(\Lab_UT.scdp.N_378_cascade_ ));
    InMux I__3682 (
            .O(N__17310),
            .I(N__17307));
    LocalMux I__3681 (
            .O(N__17307),
            .I(N__17303));
    InMux I__3680 (
            .O(N__17306),
            .I(N__17300));
    Span4Mux_h I__3679 (
            .O(N__17303),
            .I(N__17297));
    LocalMux I__3678 (
            .O(N__17300),
            .I(\Lab_UT.scdp.byteToDecrypt_4 ));
    Odrv4 I__3677 (
            .O(N__17297),
            .I(\Lab_UT.scdp.byteToDecrypt_4 ));
    InMux I__3676 (
            .O(N__17292),
            .I(N__17288));
    InMux I__3675 (
            .O(N__17291),
            .I(N__17285));
    LocalMux I__3674 (
            .O(N__17288),
            .I(\Lab_UT.scdp.val_i_0_0 ));
    LocalMux I__3673 (
            .O(N__17285),
            .I(\Lab_UT.scdp.val_i_0_0 ));
    CascadeMux I__3672 (
            .O(N__17280),
            .I(N__17277));
    InMux I__3671 (
            .O(N__17277),
            .I(N__17271));
    InMux I__3670 (
            .O(N__17276),
            .I(N__17271));
    LocalMux I__3669 (
            .O(N__17271),
            .I(\Lab_UT.scdp.N_378 ));
    CascadeMux I__3668 (
            .O(N__17268),
            .I(N__17264));
    InMux I__3667 (
            .O(N__17267),
            .I(N__17259));
    InMux I__3666 (
            .O(N__17264),
            .I(N__17252));
    InMux I__3665 (
            .O(N__17263),
            .I(N__17252));
    InMux I__3664 (
            .O(N__17262),
            .I(N__17252));
    LocalMux I__3663 (
            .O(N__17259),
            .I(N__17248));
    LocalMux I__3662 (
            .O(N__17252),
            .I(N__17245));
    InMux I__3661 (
            .O(N__17251),
            .I(N__17242));
    Span4Mux_h I__3660 (
            .O(N__17248),
            .I(N__17237));
    Span4Mux_v I__3659 (
            .O(N__17245),
            .I(N__17237));
    LocalMux I__3658 (
            .O(N__17242),
            .I(\Lab_UT.scdp.u1.byteToDecryptZ0Z_0 ));
    Odrv4 I__3657 (
            .O(N__17237),
            .I(\Lab_UT.scdp.u1.byteToDecryptZ0Z_0 ));
    InMux I__3656 (
            .O(N__17232),
            .I(N__17229));
    LocalMux I__3655 (
            .O(N__17229),
            .I(N__17226));
    Span4Mux_v I__3654 (
            .O(N__17226),
            .I(N__17223));
    Span4Mux_h I__3653 (
            .O(N__17223),
            .I(N__17220));
    Odrv4 I__3652 (
            .O(N__17220),
            .I(\Lab_UT.scdp.a2b.val_0_tz_0_3 ));
    CascadeMux I__3651 (
            .O(N__17217),
            .I(N__17214));
    InMux I__3650 (
            .O(N__17214),
            .I(N__17207));
    InMux I__3649 (
            .O(N__17213),
            .I(N__17207));
    InMux I__3648 (
            .O(N__17212),
            .I(N__17202));
    LocalMux I__3647 (
            .O(N__17207),
            .I(N__17199));
    CascadeMux I__3646 (
            .O(N__17206),
            .I(N__17192));
    InMux I__3645 (
            .O(N__17205),
            .I(N__17187));
    LocalMux I__3644 (
            .O(N__17202),
            .I(N__17182));
    Span4Mux_s3_v I__3643 (
            .O(N__17199),
            .I(N__17182));
    InMux I__3642 (
            .O(N__17198),
            .I(N__17175));
    InMux I__3641 (
            .O(N__17197),
            .I(N__17175));
    InMux I__3640 (
            .O(N__17196),
            .I(N__17175));
    InMux I__3639 (
            .O(N__17195),
            .I(N__17172));
    InMux I__3638 (
            .O(N__17192),
            .I(N__17167));
    InMux I__3637 (
            .O(N__17191),
            .I(N__17167));
    CascadeMux I__3636 (
            .O(N__17190),
            .I(N__17156));
    LocalMux I__3635 (
            .O(N__17187),
            .I(N__17152));
    Span4Mux_v I__3634 (
            .O(N__17182),
            .I(N__17147));
    LocalMux I__3633 (
            .O(N__17175),
            .I(N__17147));
    LocalMux I__3632 (
            .O(N__17172),
            .I(N__17142));
    LocalMux I__3631 (
            .O(N__17167),
            .I(N__17142));
    InMux I__3630 (
            .O(N__17166),
            .I(N__17133));
    InMux I__3629 (
            .O(N__17165),
            .I(N__17133));
    InMux I__3628 (
            .O(N__17164),
            .I(N__17133));
    InMux I__3627 (
            .O(N__17163),
            .I(N__17133));
    InMux I__3626 (
            .O(N__17162),
            .I(N__17130));
    InMux I__3625 (
            .O(N__17161),
            .I(N__17125));
    InMux I__3624 (
            .O(N__17160),
            .I(N__17118));
    InMux I__3623 (
            .O(N__17159),
            .I(N__17118));
    InMux I__3622 (
            .O(N__17156),
            .I(N__17118));
    InMux I__3621 (
            .O(N__17155),
            .I(N__17115));
    Span4Mux_v I__3620 (
            .O(N__17152),
            .I(N__17110));
    Span4Mux_v I__3619 (
            .O(N__17147),
            .I(N__17110));
    Span4Mux_v I__3618 (
            .O(N__17142),
            .I(N__17107));
    LocalMux I__3617 (
            .O(N__17133),
            .I(N__17102));
    LocalMux I__3616 (
            .O(N__17130),
            .I(N__17102));
    InMux I__3615 (
            .O(N__17129),
            .I(N__17099));
    InMux I__3614 (
            .O(N__17128),
            .I(N__17096));
    LocalMux I__3613 (
            .O(N__17125),
            .I(N__17091));
    LocalMux I__3612 (
            .O(N__17118),
            .I(N__17091));
    LocalMux I__3611 (
            .O(N__17115),
            .I(bu_rx_data_1));
    Odrv4 I__3610 (
            .O(N__17110),
            .I(bu_rx_data_1));
    Odrv4 I__3609 (
            .O(N__17107),
            .I(bu_rx_data_1));
    Odrv12 I__3608 (
            .O(N__17102),
            .I(bu_rx_data_1));
    LocalMux I__3607 (
            .O(N__17099),
            .I(bu_rx_data_1));
    LocalMux I__3606 (
            .O(N__17096),
            .I(bu_rx_data_1));
    Odrv4 I__3605 (
            .O(N__17091),
            .I(bu_rx_data_1));
    CascadeMux I__3604 (
            .O(N__17076),
            .I(N__17071));
    InMux I__3603 (
            .O(N__17075),
            .I(N__17064));
    InMux I__3602 (
            .O(N__17074),
            .I(N__17064));
    InMux I__3601 (
            .O(N__17071),
            .I(N__17064));
    LocalMux I__3600 (
            .O(N__17064),
            .I(N__17061));
    Span4Mux_v I__3599 (
            .O(N__17061),
            .I(N__17058));
    Odrv4 I__3598 (
            .O(N__17058),
            .I(bu_rx_data_i_2_2));
    InMux I__3597 (
            .O(N__17055),
            .I(N__17044));
    InMux I__3596 (
            .O(N__17054),
            .I(N__17044));
    CascadeMux I__3595 (
            .O(N__17053),
            .I(N__17038));
    InMux I__3594 (
            .O(N__17052),
            .I(N__17027));
    InMux I__3593 (
            .O(N__17051),
            .I(N__17027));
    InMux I__3592 (
            .O(N__17050),
            .I(N__17027));
    InMux I__3591 (
            .O(N__17049),
            .I(N__17027));
    LocalMux I__3590 (
            .O(N__17044),
            .I(N__17024));
    InMux I__3589 (
            .O(N__17043),
            .I(N__17019));
    InMux I__3588 (
            .O(N__17042),
            .I(N__17008));
    InMux I__3587 (
            .O(N__17041),
            .I(N__17008));
    InMux I__3586 (
            .O(N__17038),
            .I(N__17008));
    InMux I__3585 (
            .O(N__17037),
            .I(N__17008));
    InMux I__3584 (
            .O(N__17036),
            .I(N__17008));
    LocalMux I__3583 (
            .O(N__17027),
            .I(N__17005));
    Span4Mux_v I__3582 (
            .O(N__17024),
            .I(N__17002));
    InMux I__3581 (
            .O(N__17023),
            .I(N__16997));
    InMux I__3580 (
            .O(N__17022),
            .I(N__16997));
    LocalMux I__3579 (
            .O(N__17019),
            .I(N__16992));
    LocalMux I__3578 (
            .O(N__17008),
            .I(N__16992));
    Span4Mux_v I__3577 (
            .O(N__17005),
            .I(N__16983));
    Span4Mux_h I__3576 (
            .O(N__17002),
            .I(N__16983));
    LocalMux I__3575 (
            .O(N__16997),
            .I(N__16980));
    Span4Mux_v I__3574 (
            .O(N__16992),
            .I(N__16977));
    InMux I__3573 (
            .O(N__16991),
            .I(N__16972));
    InMux I__3572 (
            .O(N__16990),
            .I(N__16972));
    InMux I__3571 (
            .O(N__16989),
            .I(N__16967));
    InMux I__3570 (
            .O(N__16988),
            .I(N__16967));
    Odrv4 I__3569 (
            .O(N__16983),
            .I(bu_rx_data_i_2_0));
    Odrv4 I__3568 (
            .O(N__16980),
            .I(bu_rx_data_i_2_0));
    Odrv4 I__3567 (
            .O(N__16977),
            .I(bu_rx_data_i_2_0));
    LocalMux I__3566 (
            .O(N__16972),
            .I(bu_rx_data_i_2_0));
    LocalMux I__3565 (
            .O(N__16967),
            .I(bu_rx_data_i_2_0));
    InMux I__3564 (
            .O(N__16956),
            .I(N__16953));
    LocalMux I__3563 (
            .O(N__16953),
            .I(N__16948));
    InMux I__3562 (
            .O(N__16952),
            .I(N__16943));
    InMux I__3561 (
            .O(N__16951),
            .I(N__16943));
    Span4Mux_v I__3560 (
            .O(N__16948),
            .I(N__16940));
    LocalMux I__3559 (
            .O(N__16943),
            .I(N__16937));
    Odrv4 I__3558 (
            .O(N__16940),
            .I(\Lab_UT.sccDnibble1En ));
    Odrv4 I__3557 (
            .O(N__16937),
            .I(\Lab_UT.sccDnibble1En ));
    CascadeMux I__3556 (
            .O(N__16932),
            .I(\Lab_UT.scdp.val_0_tz_3_cascade_ ));
    InMux I__3555 (
            .O(N__16929),
            .I(N__16919));
    InMux I__3554 (
            .O(N__16928),
            .I(N__16919));
    InMux I__3553 (
            .O(N__16927),
            .I(N__16919));
    InMux I__3552 (
            .O(N__16926),
            .I(N__16916));
    LocalMux I__3551 (
            .O(N__16919),
            .I(N__16913));
    LocalMux I__3550 (
            .O(N__16916),
            .I(\Lab_UT.scdp.byteToDecrypt_7 ));
    Odrv12 I__3549 (
            .O(N__16913),
            .I(\Lab_UT.scdp.byteToDecrypt_7 ));
    InMux I__3548 (
            .O(N__16908),
            .I(N__16904));
    CascadeMux I__3547 (
            .O(N__16907),
            .I(N__16901));
    LocalMux I__3546 (
            .O(N__16904),
            .I(N__16898));
    InMux I__3545 (
            .O(N__16901),
            .I(N__16895));
    Odrv12 I__3544 (
            .O(N__16898),
            .I(\Lab_UT.scdp.key2_0 ));
    LocalMux I__3543 (
            .O(N__16895),
            .I(\Lab_UT.scdp.key2_0 ));
    InMux I__3542 (
            .O(N__16890),
            .I(N__16887));
    LocalMux I__3541 (
            .O(N__16887),
            .I(N__16883));
    CascadeMux I__3540 (
            .O(N__16886),
            .I(N__16880));
    Span12Mux_s3_v I__3539 (
            .O(N__16883),
            .I(N__16877));
    InMux I__3538 (
            .O(N__16880),
            .I(N__16874));
    Odrv12 I__3537 (
            .O(N__16877),
            .I(\Lab_UT.scdp.key2_1 ));
    LocalMux I__3536 (
            .O(N__16874),
            .I(\Lab_UT.scdp.key2_1 ));
    InMux I__3535 (
            .O(N__16869),
            .I(N__16865));
    CascadeMux I__3534 (
            .O(N__16868),
            .I(N__16862));
    LocalMux I__3533 (
            .O(N__16865),
            .I(N__16859));
    InMux I__3532 (
            .O(N__16862),
            .I(N__16856));
    Odrv4 I__3531 (
            .O(N__16859),
            .I(\Lab_UT.scdp.key3_0 ));
    LocalMux I__3530 (
            .O(N__16856),
            .I(\Lab_UT.scdp.key3_0 ));
    InMux I__3529 (
            .O(N__16851),
            .I(N__16848));
    LocalMux I__3528 (
            .O(N__16848),
            .I(N__16845));
    Span4Mux_h I__3527 (
            .O(N__16845),
            .I(N__16841));
    CascadeMux I__3526 (
            .O(N__16844),
            .I(N__16838));
    Span4Mux_h I__3525 (
            .O(N__16841),
            .I(N__16835));
    InMux I__3524 (
            .O(N__16838),
            .I(N__16832));
    Odrv4 I__3523 (
            .O(N__16835),
            .I(\Lab_UT.scdp.key3_1 ));
    LocalMux I__3522 (
            .O(N__16832),
            .I(\Lab_UT.scdp.key3_1 ));
    CascadeMux I__3521 (
            .O(N__16827),
            .I(N__16821));
    InMux I__3520 (
            .O(N__16826),
            .I(N__16817));
    InMux I__3519 (
            .O(N__16825),
            .I(N__16808));
    InMux I__3518 (
            .O(N__16824),
            .I(N__16808));
    InMux I__3517 (
            .O(N__16821),
            .I(N__16808));
    InMux I__3516 (
            .O(N__16820),
            .I(N__16808));
    LocalMux I__3515 (
            .O(N__16817),
            .I(N__16805));
    LocalMux I__3514 (
            .O(N__16808),
            .I(N__16802));
    Span4Mux_h I__3513 (
            .O(N__16805),
            .I(N__16796));
    Span4Mux_v I__3512 (
            .O(N__16802),
            .I(N__16793));
    InMux I__3511 (
            .O(N__16801),
            .I(N__16790));
    InMux I__3510 (
            .O(N__16800),
            .I(N__16785));
    InMux I__3509 (
            .O(N__16799),
            .I(N__16785));
    Odrv4 I__3508 (
            .O(N__16796),
            .I(\Lab_UT.scdp.binValD_2 ));
    Odrv4 I__3507 (
            .O(N__16793),
            .I(\Lab_UT.scdp.binValD_2 ));
    LocalMux I__3506 (
            .O(N__16790),
            .I(\Lab_UT.scdp.binValD_2 ));
    LocalMux I__3505 (
            .O(N__16785),
            .I(\Lab_UT.scdp.binValD_2 ));
    InMux I__3504 (
            .O(N__16776),
            .I(N__16773));
    LocalMux I__3503 (
            .O(N__16773),
            .I(N__16769));
    CascadeMux I__3502 (
            .O(N__16772),
            .I(N__16766));
    Span4Mux_s3_v I__3501 (
            .O(N__16769),
            .I(N__16763));
    InMux I__3500 (
            .O(N__16766),
            .I(N__16760));
    Odrv4 I__3499 (
            .O(N__16763),
            .I(\Lab_UT.scdp.key3_2 ));
    LocalMux I__3498 (
            .O(N__16760),
            .I(\Lab_UT.scdp.key3_2 ));
    InMux I__3497 (
            .O(N__16755),
            .I(N__16752));
    LocalMux I__3496 (
            .O(N__16752),
            .I(N__16749));
    Span4Mux_v I__3495 (
            .O(N__16749),
            .I(N__16746));
    Odrv4 I__3494 (
            .O(N__16746),
            .I(\Lab_UT.scctrl.g1_1_0 ));
    InMux I__3493 (
            .O(N__16743),
            .I(N__16740));
    LocalMux I__3492 (
            .O(N__16740),
            .I(\Lab_UT.scctrl.N_444_1_0 ));
    InMux I__3491 (
            .O(N__16737),
            .I(N__16731));
    InMux I__3490 (
            .O(N__16736),
            .I(N__16731));
    LocalMux I__3489 (
            .O(N__16731),
            .I(N__16727));
    InMux I__3488 (
            .O(N__16730),
            .I(N__16724));
    Odrv4 I__3487 (
            .O(N__16727),
            .I(\Lab_UT.scctrl.g0_1_1 ));
    LocalMux I__3486 (
            .O(N__16724),
            .I(\Lab_UT.scctrl.g0_1_1 ));
    CascadeMux I__3485 (
            .O(N__16719),
            .I(\Lab_UT.scctrl.g1_0_3_cascade_ ));
    InMux I__3484 (
            .O(N__16716),
            .I(N__16713));
    LocalMux I__3483 (
            .O(N__16713),
            .I(\Lab_UT.scctrl.g1_2 ));
    InMux I__3482 (
            .O(N__16710),
            .I(N__16707));
    LocalMux I__3481 (
            .O(N__16707),
            .I(\Lab_UT.scctrl.N_418_0_0 ));
    CascadeMux I__3480 (
            .O(N__16704),
            .I(N__16700));
    InMux I__3479 (
            .O(N__16703),
            .I(N__16697));
    InMux I__3478 (
            .O(N__16700),
            .I(N__16694));
    LocalMux I__3477 (
            .O(N__16697),
            .I(N__16691));
    LocalMux I__3476 (
            .O(N__16694),
            .I(N__16688));
    Span4Mux_v I__3475 (
            .O(N__16691),
            .I(N__16685));
    Span4Mux_v I__3474 (
            .O(N__16688),
            .I(N__16682));
    Odrv4 I__3473 (
            .O(N__16685),
            .I(\Lab_UT.scctrl.g0_0 ));
    Odrv4 I__3472 (
            .O(N__16682),
            .I(\Lab_UT.scctrl.g0_0 ));
    InMux I__3471 (
            .O(N__16677),
            .I(N__16674));
    LocalMux I__3470 (
            .O(N__16674),
            .I(\Lab_UT.scctrl.g0_2_1 ));
    InMux I__3469 (
            .O(N__16671),
            .I(N__16668));
    LocalMux I__3468 (
            .O(N__16668),
            .I(\Lab_UT.scctrl.g0_9_a2_2 ));
    InMux I__3467 (
            .O(N__16665),
            .I(N__16662));
    LocalMux I__3466 (
            .O(N__16662),
            .I(N__16658));
    InMux I__3465 (
            .O(N__16661),
            .I(N__16655));
    Span12Mux_s4_v I__3464 (
            .O(N__16658),
            .I(N__16652));
    LocalMux I__3463 (
            .O(N__16655),
            .I(\Lab_UT.scdp.byteToDecrypt_3 ));
    Odrv12 I__3462 (
            .O(N__16652),
            .I(\Lab_UT.scdp.byteToDecrypt_3 ));
    CascadeMux I__3461 (
            .O(N__16647),
            .I(\Lab_UT.scdp.val_i_0_0_cascade_ ));
    InMux I__3460 (
            .O(N__16644),
            .I(N__16635));
    InMux I__3459 (
            .O(N__16643),
            .I(N__16632));
    InMux I__3458 (
            .O(N__16642),
            .I(N__16629));
    CascadeMux I__3457 (
            .O(N__16641),
            .I(N__16626));
    CascadeMux I__3456 (
            .O(N__16640),
            .I(N__16623));
    CascadeMux I__3455 (
            .O(N__16639),
            .I(N__16620));
    CascadeMux I__3454 (
            .O(N__16638),
            .I(N__16617));
    LocalMux I__3453 (
            .O(N__16635),
            .I(N__16612));
    LocalMux I__3452 (
            .O(N__16632),
            .I(N__16612));
    LocalMux I__3451 (
            .O(N__16629),
            .I(N__16609));
    InMux I__3450 (
            .O(N__16626),
            .I(N__16604));
    InMux I__3449 (
            .O(N__16623),
            .I(N__16604));
    InMux I__3448 (
            .O(N__16620),
            .I(N__16599));
    InMux I__3447 (
            .O(N__16617),
            .I(N__16599));
    Span4Mux_v I__3446 (
            .O(N__16612),
            .I(N__16596));
    Span4Mux_v I__3445 (
            .O(N__16609),
            .I(N__16589));
    LocalMux I__3444 (
            .O(N__16604),
            .I(N__16589));
    LocalMux I__3443 (
            .O(N__16599),
            .I(N__16589));
    Span4Mux_v I__3442 (
            .O(N__16596),
            .I(N__16584));
    Span4Mux_v I__3441 (
            .O(N__16589),
            .I(N__16584));
    Odrv4 I__3440 (
            .O(N__16584),
            .I(\Lab_UT.scdp.a2b.N_280 ));
    CascadeMux I__3439 (
            .O(N__16581),
            .I(N__16577));
    InMux I__3438 (
            .O(N__16580),
            .I(N__16572));
    InMux I__3437 (
            .O(N__16577),
            .I(N__16569));
    InMux I__3436 (
            .O(N__16576),
            .I(N__16566));
    CascadeMux I__3435 (
            .O(N__16575),
            .I(N__16563));
    LocalMux I__3434 (
            .O(N__16572),
            .I(N__16556));
    LocalMux I__3433 (
            .O(N__16569),
            .I(N__16553));
    LocalMux I__3432 (
            .O(N__16566),
            .I(N__16550));
    InMux I__3431 (
            .O(N__16563),
            .I(N__16547));
    InMux I__3430 (
            .O(N__16562),
            .I(N__16544));
    InMux I__3429 (
            .O(N__16561),
            .I(N__16539));
    InMux I__3428 (
            .O(N__16560),
            .I(N__16539));
    InMux I__3427 (
            .O(N__16559),
            .I(N__16536));
    Span4Mux_v I__3426 (
            .O(N__16556),
            .I(N__16533));
    Span4Mux_v I__3425 (
            .O(N__16553),
            .I(N__16530));
    Span4Mux_h I__3424 (
            .O(N__16550),
            .I(N__16527));
    LocalMux I__3423 (
            .O(N__16547),
            .I(N__16524));
    LocalMux I__3422 (
            .O(N__16544),
            .I(N__16521));
    LocalMux I__3421 (
            .O(N__16539),
            .I(N__16516));
    LocalMux I__3420 (
            .O(N__16536),
            .I(N__16516));
    Span4Mux_h I__3419 (
            .O(N__16533),
            .I(N__16507));
    Span4Mux_s2_h I__3418 (
            .O(N__16530),
            .I(N__16507));
    Span4Mux_v I__3417 (
            .O(N__16527),
            .I(N__16507));
    Span4Mux_v I__3416 (
            .O(N__16524),
            .I(N__16507));
    Span4Mux_v I__3415 (
            .O(N__16521),
            .I(N__16502));
    Span4Mux_v I__3414 (
            .O(N__16516),
            .I(N__16502));
    Odrv4 I__3413 (
            .O(N__16507),
            .I(bu_rx_data_0));
    Odrv4 I__3412 (
            .O(N__16502),
            .I(bu_rx_data_0));
    CEMux I__3411 (
            .O(N__16497),
            .I(N__16494));
    LocalMux I__3410 (
            .O(N__16494),
            .I(N__16491));
    Span4Mux_v I__3409 (
            .O(N__16491),
            .I(N__16488));
    Odrv4 I__3408 (
            .O(N__16488),
            .I(\Lab_UT.scctrl.N_398i_i ));
    CascadeMux I__3407 (
            .O(N__16485),
            .I(N__16482));
    InMux I__3406 (
            .O(N__16482),
            .I(N__16479));
    LocalMux I__3405 (
            .O(N__16479),
            .I(N__16476));
    Span4Mux_v I__3404 (
            .O(N__16476),
            .I(N__16473));
    Span4Mux_h I__3403 (
            .O(N__16473),
            .I(N__16470));
    Odrv4 I__3402 (
            .O(N__16470),
            .I(\Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0_0 ));
    InMux I__3401 (
            .O(N__16467),
            .I(N__16461));
    InMux I__3400 (
            .O(N__16466),
            .I(N__16461));
    LocalMux I__3399 (
            .O(N__16461),
            .I(\Lab_UT.scctrl.nibbleInZ0Z1 ));
    CascadeMux I__3398 (
            .O(N__16458),
            .I(\Lab_UT.scctrl.N_69_cascade_ ));
    CascadeMux I__3397 (
            .O(N__16455),
            .I(\Lab_UT.sccDnibble1En_cascade_ ));
    InMux I__3396 (
            .O(N__16452),
            .I(N__16448));
    IoInMux I__3395 (
            .O(N__16451),
            .I(N__16444));
    LocalMux I__3394 (
            .O(N__16448),
            .I(N__16441));
    InMux I__3393 (
            .O(N__16447),
            .I(N__16438));
    LocalMux I__3392 (
            .O(N__16444),
            .I(N__16435));
    Span4Mux_h I__3391 (
            .O(N__16441),
            .I(N__16432));
    LocalMux I__3390 (
            .O(N__16438),
            .I(N__16429));
    IoSpan4Mux I__3389 (
            .O(N__16435),
            .I(N__16426));
    Span4Mux_h I__3388 (
            .O(N__16432),
            .I(N__16423));
    Span4Mux_v I__3387 (
            .O(N__16429),
            .I(N__16420));
    Span4Mux_s3_h I__3386 (
            .O(N__16426),
            .I(N__16417));
    Odrv4 I__3385 (
            .O(N__16423),
            .I(resetGen_rst_1_iso));
    Odrv4 I__3384 (
            .O(N__16420),
            .I(resetGen_rst_1_iso));
    Odrv4 I__3383 (
            .O(N__16417),
            .I(resetGen_rst_1_iso));
    CEMux I__3382 (
            .O(N__16410),
            .I(N__16407));
    LocalMux I__3381 (
            .O(N__16407),
            .I(N__16404));
    Span4Mux_h I__3380 (
            .O(N__16404),
            .I(N__16401));
    Span4Mux_v I__3379 (
            .O(N__16401),
            .I(N__16398));
    Odrv4 I__3378 (
            .O(N__16398),
            .I(\Lab_UT.scdp.u0.sccDnibble1En_0 ));
    InMux I__3377 (
            .O(N__16395),
            .I(N__16392));
    LocalMux I__3376 (
            .O(N__16392),
            .I(N__16389));
    Span4Mux_s3_h I__3375 (
            .O(N__16389),
            .I(N__16386));
    Span4Mux_h I__3374 (
            .O(N__16386),
            .I(N__16383));
    Odrv4 I__3373 (
            .O(N__16383),
            .I(\Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0dup_1 ));
    InMux I__3372 (
            .O(N__16380),
            .I(N__16377));
    LocalMux I__3371 (
            .O(N__16377),
            .I(\Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93 ));
    CascadeMux I__3370 (
            .O(N__16374),
            .I(\Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93_cascade_ ));
    SRMux I__3369 (
            .O(N__16371),
            .I(N__16368));
    LocalMux I__3368 (
            .O(N__16368),
            .I(\Lab_UT.scctrl.N_69_i ));
    InMux I__3367 (
            .O(N__16365),
            .I(N__16362));
    LocalMux I__3366 (
            .O(N__16362),
            .I(\Lab_UT.scctrl.N_11 ));
    CascadeMux I__3365 (
            .O(N__16359),
            .I(N__16355));
    InMux I__3364 (
            .O(N__16358),
            .I(N__16349));
    InMux I__3363 (
            .O(N__16355),
            .I(N__16340));
    InMux I__3362 (
            .O(N__16354),
            .I(N__16340));
    InMux I__3361 (
            .O(N__16353),
            .I(N__16340));
    InMux I__3360 (
            .O(N__16352),
            .I(N__16340));
    LocalMux I__3359 (
            .O(N__16349),
            .I(N__16337));
    LocalMux I__3358 (
            .O(N__16340),
            .I(\Lab_UT.scctrl.next_state_rst ));
    Odrv4 I__3357 (
            .O(N__16337),
            .I(\Lab_UT.scctrl.next_state_rst ));
    CascadeMux I__3356 (
            .O(N__16332),
            .I(\Lab_UT.scctrl.g0_9_a2_5_cascade_ ));
    InMux I__3355 (
            .O(N__16329),
            .I(N__16323));
    InMux I__3354 (
            .O(N__16328),
            .I(N__16323));
    LocalMux I__3353 (
            .O(N__16323),
            .I(\Lab_UT.scctrl.next_state_rst_0_3_tz ));
    CascadeMux I__3352 (
            .O(N__16320),
            .I(\Lab_UT.scctrl.next_state_rst_0_3_0_cascade_ ));
    InMux I__3351 (
            .O(N__16317),
            .I(N__16313));
    CascadeMux I__3350 (
            .O(N__16316),
            .I(N__16310));
    LocalMux I__3349 (
            .O(N__16313),
            .I(N__16307));
    InMux I__3348 (
            .O(N__16310),
            .I(N__16302));
    Span4Mux_v I__3347 (
            .O(N__16307),
            .I(N__16299));
    InMux I__3346 (
            .O(N__16306),
            .I(N__16296));
    InMux I__3345 (
            .O(N__16305),
            .I(N__16293));
    LocalMux I__3344 (
            .O(N__16302),
            .I(N__16288));
    Span4Mux_s2_h I__3343 (
            .O(N__16299),
            .I(N__16288));
    LocalMux I__3342 (
            .O(N__16296),
            .I(rst_i_fast));
    LocalMux I__3341 (
            .O(N__16293),
            .I(rst_i_fast));
    Odrv4 I__3340 (
            .O(N__16288),
            .I(rst_i_fast));
    InMux I__3339 (
            .O(N__16281),
            .I(N__16276));
    InMux I__3338 (
            .O(N__16280),
            .I(N__16273));
    InMux I__3337 (
            .O(N__16279),
            .I(N__16270));
    LocalMux I__3336 (
            .O(N__16276),
            .I(N__16267));
    LocalMux I__3335 (
            .O(N__16273),
            .I(N__16264));
    LocalMux I__3334 (
            .O(N__16270),
            .I(\Lab_UT.scctrl.state_fast_3 ));
    Odrv12 I__3333 (
            .O(N__16267),
            .I(\Lab_UT.scctrl.state_fast_3 ));
    Odrv4 I__3332 (
            .O(N__16264),
            .I(\Lab_UT.scctrl.state_fast_3 ));
    CascadeMux I__3331 (
            .O(N__16257),
            .I(\Lab_UT.scctrl.g0_0_0_0_cascade_ ));
    CascadeMux I__3330 (
            .O(N__16254),
            .I(\Lab_UT.scctrl.g0_0_2_cascade_ ));
    InMux I__3329 (
            .O(N__16251),
            .I(N__16248));
    LocalMux I__3328 (
            .O(N__16248),
            .I(\Lab_UT.scctrl.g0_0_3 ));
    InMux I__3327 (
            .O(N__16245),
            .I(N__16242));
    LocalMux I__3326 (
            .O(N__16242),
            .I(N__16238));
    InMux I__3325 (
            .O(N__16241),
            .I(N__16235));
    Odrv4 I__3324 (
            .O(N__16238),
            .I(buart__rx_shifter_1_fast_0));
    LocalMux I__3323 (
            .O(N__16235),
            .I(buart__rx_shifter_1_fast_0));
    InMux I__3322 (
            .O(N__16230),
            .I(N__16227));
    LocalMux I__3321 (
            .O(N__16227),
            .I(\Lab_UT.scctrl.N_408_0 ));
    InMux I__3320 (
            .O(N__16224),
            .I(N__16221));
    LocalMux I__3319 (
            .O(N__16221),
            .I(\Lab_UT.scctrl.g2_0_0 ));
    InMux I__3318 (
            .O(N__16218),
            .I(N__16215));
    LocalMux I__3317 (
            .O(N__16215),
            .I(\Lab_UT.scctrl.N_17 ));
    InMux I__3316 (
            .O(N__16212),
            .I(N__16201));
    InMux I__3315 (
            .O(N__16211),
            .I(N__16201));
    InMux I__3314 (
            .O(N__16210),
            .I(N__16198));
    InMux I__3313 (
            .O(N__16209),
            .I(N__16193));
    InMux I__3312 (
            .O(N__16208),
            .I(N__16193));
    InMux I__3311 (
            .O(N__16207),
            .I(N__16186));
    InMux I__3310 (
            .O(N__16206),
            .I(N__16186));
    LocalMux I__3309 (
            .O(N__16201),
            .I(N__16183));
    LocalMux I__3308 (
            .O(N__16198),
            .I(N__16178));
    LocalMux I__3307 (
            .O(N__16193),
            .I(N__16178));
    InMux I__3306 (
            .O(N__16192),
            .I(N__16173));
    InMux I__3305 (
            .O(N__16191),
            .I(N__16173));
    LocalMux I__3304 (
            .O(N__16186),
            .I(\Lab_UT.scctrl.N_240_i_0 ));
    Odrv4 I__3303 (
            .O(N__16183),
            .I(\Lab_UT.scctrl.N_240_i_0 ));
    Odrv12 I__3302 (
            .O(N__16178),
            .I(\Lab_UT.scctrl.N_240_i_0 ));
    LocalMux I__3301 (
            .O(N__16173),
            .I(\Lab_UT.scctrl.N_240_i_0 ));
    CascadeMux I__3300 (
            .O(N__16164),
            .I(N__16159));
    InMux I__3299 (
            .O(N__16163),
            .I(N__16139));
    InMux I__3298 (
            .O(N__16162),
            .I(N__16139));
    InMux I__3297 (
            .O(N__16159),
            .I(N__16139));
    InMux I__3296 (
            .O(N__16158),
            .I(N__16135));
    InMux I__3295 (
            .O(N__16157),
            .I(N__16132));
    InMux I__3294 (
            .O(N__16156),
            .I(N__16121));
    InMux I__3293 (
            .O(N__16155),
            .I(N__16121));
    InMux I__3292 (
            .O(N__16154),
            .I(N__16121));
    InMux I__3291 (
            .O(N__16153),
            .I(N__16121));
    InMux I__3290 (
            .O(N__16152),
            .I(N__16121));
    InMux I__3289 (
            .O(N__16151),
            .I(N__16118));
    InMux I__3288 (
            .O(N__16150),
            .I(N__16113));
    InMux I__3287 (
            .O(N__16149),
            .I(N__16113));
    InMux I__3286 (
            .O(N__16148),
            .I(N__16108));
    InMux I__3285 (
            .O(N__16147),
            .I(N__16108));
    CascadeMux I__3284 (
            .O(N__16146),
            .I(N__16105));
    LocalMux I__3283 (
            .O(N__16139),
            .I(N__16101));
    InMux I__3282 (
            .O(N__16138),
            .I(N__16096));
    LocalMux I__3281 (
            .O(N__16135),
            .I(N__16093));
    LocalMux I__3280 (
            .O(N__16132),
            .I(N__16088));
    LocalMux I__3279 (
            .O(N__16121),
            .I(N__16088));
    LocalMux I__3278 (
            .O(N__16118),
            .I(N__16081));
    LocalMux I__3277 (
            .O(N__16113),
            .I(N__16081));
    LocalMux I__3276 (
            .O(N__16108),
            .I(N__16081));
    InMux I__3275 (
            .O(N__16105),
            .I(N__16078));
    InMux I__3274 (
            .O(N__16104),
            .I(N__16075));
    Span4Mux_v I__3273 (
            .O(N__16101),
            .I(N__16072));
    InMux I__3272 (
            .O(N__16100),
            .I(N__16067));
    InMux I__3271 (
            .O(N__16099),
            .I(N__16067));
    LocalMux I__3270 (
            .O(N__16096),
            .I(N__16056));
    Span4Mux_v I__3269 (
            .O(N__16093),
            .I(N__16056));
    Span4Mux_v I__3268 (
            .O(N__16088),
            .I(N__16056));
    Span4Mux_v I__3267 (
            .O(N__16081),
            .I(N__16056));
    LocalMux I__3266 (
            .O(N__16078),
            .I(N__16056));
    LocalMux I__3265 (
            .O(N__16075),
            .I(N__16051));
    Span4Mux_s2_h I__3264 (
            .O(N__16072),
            .I(N__16051));
    LocalMux I__3263 (
            .O(N__16067),
            .I(bu_rx_data_i_1_5));
    Odrv4 I__3262 (
            .O(N__16056),
            .I(bu_rx_data_i_1_5));
    Odrv4 I__3261 (
            .O(N__16051),
            .I(bu_rx_data_i_1_5));
    CascadeMux I__3260 (
            .O(N__16044),
            .I(\Lab_UT.scctrl.N_412_cascade_ ));
    InMux I__3259 (
            .O(N__16041),
            .I(N__16035));
    InMux I__3258 (
            .O(N__16040),
            .I(N__16035));
    LocalMux I__3257 (
            .O(N__16035),
            .I(\Lab_UT.scctrl.next_state_rst_0_1 ));
    CascadeMux I__3256 (
            .O(N__16032),
            .I(\Lab_UT.scctrl.state_ret_4_RNOZ0Z_10_cascade_ ));
    InMux I__3255 (
            .O(N__16029),
            .I(N__16026));
    LocalMux I__3254 (
            .O(N__16026),
            .I(N__16023));
    Span4Mux_v I__3253 (
            .O(N__16023),
            .I(N__16020));
    Odrv4 I__3252 (
            .O(N__16020),
            .I(\Lab_UT.scctrl.state_ret_4_RNOZ0Z_6 ));
    CascadeMux I__3251 (
            .O(N__16017),
            .I(N__16014));
    InMux I__3250 (
            .O(N__16014),
            .I(N__16007));
    InMux I__3249 (
            .O(N__16013),
            .I(N__16007));
    InMux I__3248 (
            .O(N__16012),
            .I(N__16004));
    LocalMux I__3247 (
            .O(N__16007),
            .I(N__15999));
    LocalMux I__3246 (
            .O(N__16004),
            .I(N__15999));
    Span4Mux_v I__3245 (
            .O(N__15999),
            .I(N__15996));
    Odrv4 I__3244 (
            .O(N__15996),
            .I(\Lab_UT.scctrl.N_295 ));
    CascadeMux I__3243 (
            .O(N__15993),
            .I(\Lab_UT.scctrl.N_295_cascade_ ));
    InMux I__3242 (
            .O(N__15990),
            .I(N__15987));
    LocalMux I__3241 (
            .O(N__15987),
            .I(N__15984));
    Sp12to4 I__3240 (
            .O(N__15984),
            .I(N__15981));
    Odrv12 I__3239 (
            .O(N__15981),
            .I(\Lab_UT.scctrl.N_40_i ));
    InMux I__3238 (
            .O(N__15978),
            .I(N__15971));
    CascadeMux I__3237 (
            .O(N__15977),
            .I(N__15968));
    CascadeMux I__3236 (
            .O(N__15976),
            .I(N__15965));
    CascadeMux I__3235 (
            .O(N__15975),
            .I(N__15962));
    CascadeMux I__3234 (
            .O(N__15974),
            .I(N__15959));
    LocalMux I__3233 (
            .O(N__15971),
            .I(N__15956));
    InMux I__3232 (
            .O(N__15968),
            .I(N__15953));
    InMux I__3231 (
            .O(N__15965),
            .I(N__15949));
    InMux I__3230 (
            .O(N__15962),
            .I(N__15944));
    InMux I__3229 (
            .O(N__15959),
            .I(N__15944));
    Span4Mux_h I__3228 (
            .O(N__15956),
            .I(N__15941));
    LocalMux I__3227 (
            .O(N__15953),
            .I(N__15938));
    InMux I__3226 (
            .O(N__15952),
            .I(N__15935));
    LocalMux I__3225 (
            .O(N__15949),
            .I(\Lab_UT.scctrl.N_487 ));
    LocalMux I__3224 (
            .O(N__15944),
            .I(\Lab_UT.scctrl.N_487 ));
    Odrv4 I__3223 (
            .O(N__15941),
            .I(\Lab_UT.scctrl.N_487 ));
    Odrv4 I__3222 (
            .O(N__15938),
            .I(\Lab_UT.scctrl.N_487 ));
    LocalMux I__3221 (
            .O(N__15935),
            .I(\Lab_UT.scctrl.N_487 ));
    InMux I__3220 (
            .O(N__15924),
            .I(N__15921));
    LocalMux I__3219 (
            .O(N__15921),
            .I(N__15916));
    InMux I__3218 (
            .O(N__15920),
            .I(N__15911));
    InMux I__3217 (
            .O(N__15919),
            .I(N__15911));
    Span4Mux_h I__3216 (
            .O(N__15916),
            .I(N__15908));
    LocalMux I__3215 (
            .O(N__15911),
            .I(\Lab_UT.scctrl.N_284 ));
    Odrv4 I__3214 (
            .O(N__15908),
            .I(\Lab_UT.scctrl.N_284 ));
    CascadeMux I__3213 (
            .O(N__15903),
            .I(N__15897));
    InMux I__3212 (
            .O(N__15902),
            .I(N__15893));
    InMux I__3211 (
            .O(N__15901),
            .I(N__15888));
    InMux I__3210 (
            .O(N__15900),
            .I(N__15885));
    InMux I__3209 (
            .O(N__15897),
            .I(N__15880));
    InMux I__3208 (
            .O(N__15896),
            .I(N__15880));
    LocalMux I__3207 (
            .O(N__15893),
            .I(N__15875));
    InMux I__3206 (
            .O(N__15892),
            .I(N__15870));
    InMux I__3205 (
            .O(N__15891),
            .I(N__15870));
    LocalMux I__3204 (
            .O(N__15888),
            .I(N__15865));
    LocalMux I__3203 (
            .O(N__15885),
            .I(N__15865));
    LocalMux I__3202 (
            .O(N__15880),
            .I(N__15862));
    InMux I__3201 (
            .O(N__15879),
            .I(N__15859));
    InMux I__3200 (
            .O(N__15878),
            .I(N__15856));
    Span4Mux_v I__3199 (
            .O(N__15875),
            .I(N__15853));
    LocalMux I__3198 (
            .O(N__15870),
            .I(N__15842));
    Span4Mux_v I__3197 (
            .O(N__15865),
            .I(N__15842));
    Span4Mux_v I__3196 (
            .O(N__15862),
            .I(N__15842));
    LocalMux I__3195 (
            .O(N__15859),
            .I(N__15842));
    LocalMux I__3194 (
            .O(N__15856),
            .I(N__15842));
    Odrv4 I__3193 (
            .O(N__15853),
            .I(\Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0 ));
    Odrv4 I__3192 (
            .O(N__15842),
            .I(\Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0 ));
    CascadeMux I__3191 (
            .O(N__15837),
            .I(\Lab_UT.scctrl.N_408_cascade_ ));
    CascadeMux I__3190 (
            .O(N__15834),
            .I(\Lab_UT.scctrl.g0_i_a8_0_1_cascade_ ));
    InMux I__3189 (
            .O(N__15831),
            .I(N__15828));
    LocalMux I__3188 (
            .O(N__15828),
            .I(N__15825));
    Span4Mux_h I__3187 (
            .O(N__15825),
            .I(N__15822));
    Odrv4 I__3186 (
            .O(N__15822),
            .I(\Lab_UT.scctrl.G_24_i_o7_0_0 ));
    CascadeMux I__3185 (
            .O(N__15819),
            .I(\Lab_UT.scctrl.N_12_1_cascade_ ));
    CascadeMux I__3184 (
            .O(N__15816),
            .I(N__15813));
    InMux I__3183 (
            .O(N__15813),
            .I(N__15810));
    LocalMux I__3182 (
            .O(N__15810),
            .I(\Lab_UT.scctrl.N_408 ));
    CascadeMux I__3181 (
            .O(N__15807),
            .I(\Lab_UT.scctrl.N_418_2_cascade_ ));
    InMux I__3180 (
            .O(N__15804),
            .I(N__15801));
    LocalMux I__3179 (
            .O(N__15801),
            .I(N__15798));
    Span4Mux_h I__3178 (
            .O(N__15798),
            .I(N__15795));
    Odrv4 I__3177 (
            .O(N__15795),
            .I(\Lab_UT.scctrl.g1_0 ));
    InMux I__3176 (
            .O(N__15792),
            .I(N__15784));
    InMux I__3175 (
            .O(N__15791),
            .I(N__15773));
    InMux I__3174 (
            .O(N__15790),
            .I(N__15773));
    InMux I__3173 (
            .O(N__15789),
            .I(N__15773));
    InMux I__3172 (
            .O(N__15788),
            .I(N__15773));
    InMux I__3171 (
            .O(N__15787),
            .I(N__15773));
    LocalMux I__3170 (
            .O(N__15784),
            .I(N__15770));
    LocalMux I__3169 (
            .O(N__15773),
            .I(\Lab_UT.scctrl.N_418 ));
    Odrv4 I__3168 (
            .O(N__15770),
            .I(\Lab_UT.scctrl.N_418 ));
    CascadeMux I__3167 (
            .O(N__15765),
            .I(N__15761));
    InMux I__3166 (
            .O(N__15764),
            .I(N__15756));
    InMux I__3165 (
            .O(N__15761),
            .I(N__15756));
    LocalMux I__3164 (
            .O(N__15756),
            .I(N__15753));
    Span4Mux_s3_h I__3163 (
            .O(N__15753),
            .I(N__15750));
    Odrv4 I__3162 (
            .O(N__15750),
            .I(\Lab_UT.scctrl.N_415 ));
    InMux I__3161 (
            .O(N__15747),
            .I(N__15744));
    LocalMux I__3160 (
            .O(N__15744),
            .I(N__15738));
    InMux I__3159 (
            .O(N__15743),
            .I(N__15735));
    InMux I__3158 (
            .O(N__15742),
            .I(N__15730));
    InMux I__3157 (
            .O(N__15741),
            .I(N__15730));
    Span4Mux_s2_v I__3156 (
            .O(N__15738),
            .I(N__15727));
    LocalMux I__3155 (
            .O(N__15735),
            .I(\Lab_UT.scctrl.state_ret_0_fastZ0 ));
    LocalMux I__3154 (
            .O(N__15730),
            .I(\Lab_UT.scctrl.state_ret_0_fastZ0 ));
    Odrv4 I__3153 (
            .O(N__15727),
            .I(\Lab_UT.scctrl.state_ret_0_fastZ0 ));
    CascadeMux I__3152 (
            .O(N__15720),
            .I(\Lab_UT.scctrl.next_state_rst_4_4_cascade_ ));
    InMux I__3151 (
            .O(N__15717),
            .I(N__15714));
    LocalMux I__3150 (
            .O(N__15714),
            .I(\Lab_UT.scctrl.N_290_1 ));
    CascadeMux I__3149 (
            .O(N__15711),
            .I(N__15708));
    InMux I__3148 (
            .O(N__15708),
            .I(N__15705));
    LocalMux I__3147 (
            .O(N__15705),
            .I(\Lab_UT.scctrl.g0_1_0 ));
    InMux I__3146 (
            .O(N__15702),
            .I(N__15699));
    LocalMux I__3145 (
            .O(N__15699),
            .I(N__15692));
    InMux I__3144 (
            .O(N__15698),
            .I(N__15685));
    InMux I__3143 (
            .O(N__15697),
            .I(N__15685));
    InMux I__3142 (
            .O(N__15696),
            .I(N__15685));
    InMux I__3141 (
            .O(N__15695),
            .I(N__15682));
    Span4Mux_v I__3140 (
            .O(N__15692),
            .I(N__15679));
    LocalMux I__3139 (
            .O(N__15685),
            .I(\Lab_UT.scctrl.next_state_rst_1_3 ));
    LocalMux I__3138 (
            .O(N__15682),
            .I(\Lab_UT.scctrl.next_state_rst_1_3 ));
    Odrv4 I__3137 (
            .O(N__15679),
            .I(\Lab_UT.scctrl.next_state_rst_1_3 ));
    CascadeMux I__3136 (
            .O(N__15672),
            .I(\Lab_UT.scctrl.next_state_rst_4_2_cascade_ ));
    InMux I__3135 (
            .O(N__15669),
            .I(N__15666));
    LocalMux I__3134 (
            .O(N__15666),
            .I(\Lab_UT.scctrl.N_290 ));
    InMux I__3133 (
            .O(N__15663),
            .I(N__15660));
    LocalMux I__3132 (
            .O(N__15660),
            .I(N__15657));
    Odrv4 I__3131 (
            .O(N__15657),
            .I(\Lab_UT.scctrl.next_state_0_3 ));
    InMux I__3130 (
            .O(N__15654),
            .I(N__15651));
    LocalMux I__3129 (
            .O(N__15651),
            .I(\Lab_UT.scctrl.N_415_2 ));
    CascadeMux I__3128 (
            .O(N__15648),
            .I(\Lab_UT.scctrl.g1_2_0_cascade_ ));
    CascadeMux I__3127 (
            .O(N__15645),
            .I(\Lab_UT.scctrl.next_stateZ0Z_2_cascade_ ));
    InMux I__3126 (
            .O(N__15642),
            .I(N__15636));
    InMux I__3125 (
            .O(N__15641),
            .I(N__15636));
    LocalMux I__3124 (
            .O(N__15636),
            .I(N__15633));
    Span4Mux_h I__3123 (
            .O(N__15633),
            .I(N__15630));
    Span4Mux_v I__3122 (
            .O(N__15630),
            .I(N__15627));
    Odrv4 I__3121 (
            .O(N__15627),
            .I(\Lab_UT.scctrl.next_state_rst_2 ));
    CascadeMux I__3120 (
            .O(N__15624),
            .I(N__15621));
    InMux I__3119 (
            .O(N__15621),
            .I(N__15617));
    InMux I__3118 (
            .O(N__15620),
            .I(N__15614));
    LocalMux I__3117 (
            .O(N__15617),
            .I(N__15608));
    LocalMux I__3116 (
            .O(N__15614),
            .I(N__15608));
    InMux I__3115 (
            .O(N__15613),
            .I(N__15605));
    Span4Mux_v I__3114 (
            .O(N__15608),
            .I(N__15602));
    LocalMux I__3113 (
            .O(N__15605),
            .I(\Lab_UT.scctrl.next_stateZ0Z_2 ));
    Odrv4 I__3112 (
            .O(N__15602),
            .I(\Lab_UT.scctrl.next_stateZ0Z_2 ));
    CascadeMux I__3111 (
            .O(N__15597),
            .I(N__15593));
    CascadeMux I__3110 (
            .O(N__15596),
            .I(N__15590));
    InMux I__3109 (
            .O(N__15593),
            .I(N__15576));
    InMux I__3108 (
            .O(N__15590),
            .I(N__15576));
    InMux I__3107 (
            .O(N__15589),
            .I(N__15576));
    InMux I__3106 (
            .O(N__15588),
            .I(N__15576));
    InMux I__3105 (
            .O(N__15587),
            .I(N__15576));
    LocalMux I__3104 (
            .O(N__15576),
            .I(N__15573));
    Odrv4 I__3103 (
            .O(N__15573),
            .I(\Lab_UT.scctrl.g1_1_1_0 ));
    InMux I__3102 (
            .O(N__15570),
            .I(N__15558));
    InMux I__3101 (
            .O(N__15569),
            .I(N__15558));
    InMux I__3100 (
            .O(N__15568),
            .I(N__15558));
    InMux I__3099 (
            .O(N__15567),
            .I(N__15558));
    LocalMux I__3098 (
            .O(N__15558),
            .I(\Lab_UT.scctrl.g1_2_0 ));
    CascadeMux I__3097 (
            .O(N__15555),
            .I(\Lab_UT.scctrl.next_state_rst_4_3_cascade_ ));
    InMux I__3096 (
            .O(N__15552),
            .I(N__15549));
    LocalMux I__3095 (
            .O(N__15549),
            .I(N__15546));
    Odrv4 I__3094 (
            .O(N__15546),
            .I(\Lab_UT.scctrl.N_290_0 ));
    InMux I__3093 (
            .O(N__15543),
            .I(N__15540));
    LocalMux I__3092 (
            .O(N__15540),
            .I(\Lab_UT.scctrl.next_state_rst_4_5 ));
    CascadeMux I__3091 (
            .O(N__15537),
            .I(\Lab_UT.scctrl.N_20_i_cascade_ ));
    InMux I__3090 (
            .O(N__15534),
            .I(N__15531));
    LocalMux I__3089 (
            .O(N__15531),
            .I(\Lab_UT.scctrl.N_277 ));
    CascadeMux I__3088 (
            .O(N__15528),
            .I(\Lab_UT.scctrl.N_277_cascade_ ));
    IoInMux I__3087 (
            .O(N__15525),
            .I(N__15522));
    LocalMux I__3086 (
            .O(N__15522),
            .I(N__15519));
    IoSpan4Mux I__3085 (
            .O(N__15519),
            .I(N__15516));
    Span4Mux_s3_h I__3084 (
            .O(N__15516),
            .I(N__15513));
    Odrv4 I__3083 (
            .O(N__15513),
            .I(N_67));
    InMux I__3082 (
            .O(N__15510),
            .I(N__15507));
    LocalMux I__3081 (
            .O(N__15507),
            .I(\Lab_UT.scctrl.N_355 ));
    InMux I__3080 (
            .O(N__15504),
            .I(N__15500));
    InMux I__3079 (
            .O(N__15503),
            .I(N__15491));
    LocalMux I__3078 (
            .O(N__15500),
            .I(N__15488));
    InMux I__3077 (
            .O(N__15499),
            .I(N__15479));
    InMux I__3076 (
            .O(N__15498),
            .I(N__15479));
    InMux I__3075 (
            .O(N__15497),
            .I(N__15479));
    InMux I__3074 (
            .O(N__15496),
            .I(N__15479));
    InMux I__3073 (
            .O(N__15495),
            .I(N__15474));
    InMux I__3072 (
            .O(N__15494),
            .I(N__15474));
    LocalMux I__3071 (
            .O(N__15491),
            .I(\Lab_UT.scctrl.N_36 ));
    Odrv4 I__3070 (
            .O(N__15488),
            .I(\Lab_UT.scctrl.N_36 ));
    LocalMux I__3069 (
            .O(N__15479),
            .I(\Lab_UT.scctrl.N_36 ));
    LocalMux I__3068 (
            .O(N__15474),
            .I(\Lab_UT.scctrl.N_36 ));
    CascadeMux I__3067 (
            .O(N__15465),
            .I(\Lab_UT.scctrl.N_27_i_cascade_ ));
    InMux I__3066 (
            .O(N__15462),
            .I(N__15452));
    InMux I__3065 (
            .O(N__15461),
            .I(N__15444));
    InMux I__3064 (
            .O(N__15460),
            .I(N__15440));
    InMux I__3063 (
            .O(N__15459),
            .I(N__15437));
    InMux I__3062 (
            .O(N__15458),
            .I(N__15434));
    InMux I__3061 (
            .O(N__15457),
            .I(N__15431));
    InMux I__3060 (
            .O(N__15456),
            .I(N__15425));
    InMux I__3059 (
            .O(N__15455),
            .I(N__15425));
    LocalMux I__3058 (
            .O(N__15452),
            .I(N__15422));
    InMux I__3057 (
            .O(N__15451),
            .I(N__15419));
    InMux I__3056 (
            .O(N__15450),
            .I(N__15416));
    InMux I__3055 (
            .O(N__15449),
            .I(N__15411));
    InMux I__3054 (
            .O(N__15448),
            .I(N__15411));
    InMux I__3053 (
            .O(N__15447),
            .I(N__15408));
    LocalMux I__3052 (
            .O(N__15444),
            .I(N__15405));
    InMux I__3051 (
            .O(N__15443),
            .I(N__15402));
    LocalMux I__3050 (
            .O(N__15440),
            .I(N__15399));
    LocalMux I__3049 (
            .O(N__15437),
            .I(N__15395));
    LocalMux I__3048 (
            .O(N__15434),
            .I(N__15390));
    LocalMux I__3047 (
            .O(N__15431),
            .I(N__15390));
    CascadeMux I__3046 (
            .O(N__15430),
            .I(N__15387));
    LocalMux I__3045 (
            .O(N__15425),
            .I(N__15380));
    Span4Mux_h I__3044 (
            .O(N__15422),
            .I(N__15380));
    LocalMux I__3043 (
            .O(N__15419),
            .I(N__15380));
    LocalMux I__3042 (
            .O(N__15416),
            .I(N__15377));
    LocalMux I__3041 (
            .O(N__15411),
            .I(N__15374));
    LocalMux I__3040 (
            .O(N__15408),
            .I(N__15367));
    Span4Mux_v I__3039 (
            .O(N__15405),
            .I(N__15367));
    LocalMux I__3038 (
            .O(N__15402),
            .I(N__15367));
    Span4Mux_h I__3037 (
            .O(N__15399),
            .I(N__15364));
    InMux I__3036 (
            .O(N__15398),
            .I(N__15361));
    Span4Mux_v I__3035 (
            .O(N__15395),
            .I(N__15358));
    Span4Mux_h I__3034 (
            .O(N__15390),
            .I(N__15355));
    InMux I__3033 (
            .O(N__15387),
            .I(N__15352));
    Span4Mux_v I__3032 (
            .O(N__15380),
            .I(N__15347));
    Span4Mux_v I__3031 (
            .O(N__15377),
            .I(N__15347));
    Span4Mux_s3_h I__3030 (
            .O(N__15374),
            .I(N__15340));
    Span4Mux_h I__3029 (
            .O(N__15367),
            .I(N__15340));
    Span4Mux_v I__3028 (
            .O(N__15364),
            .I(N__15340));
    LocalMux I__3027 (
            .O(N__15361),
            .I(rst_i));
    Odrv4 I__3026 (
            .O(N__15358),
            .I(rst_i));
    Odrv4 I__3025 (
            .O(N__15355),
            .I(rst_i));
    LocalMux I__3024 (
            .O(N__15352),
            .I(rst_i));
    Odrv4 I__3023 (
            .O(N__15347),
            .I(rst_i));
    Odrv4 I__3022 (
            .O(N__15340),
            .I(rst_i));
    CascadeMux I__3021 (
            .O(N__15327),
            .I(N__15324));
    InMux I__3020 (
            .O(N__15324),
            .I(N__15321));
    LocalMux I__3019 (
            .O(N__15321),
            .I(\Lab_UT.scctrl.N_19 ));
    InMux I__3018 (
            .O(N__15318),
            .I(N__15315));
    LocalMux I__3017 (
            .O(N__15315),
            .I(\Lab_UT.scctrl.G_24_i_1_0 ));
    InMux I__3016 (
            .O(N__15312),
            .I(N__15308));
    InMux I__3015 (
            .O(N__15311),
            .I(N__15305));
    LocalMux I__3014 (
            .O(N__15308),
            .I(N__15302));
    LocalMux I__3013 (
            .O(N__15305),
            .I(N__15299));
    Span4Mux_h I__3012 (
            .O(N__15302),
            .I(N__15296));
    Odrv12 I__3011 (
            .O(N__15299),
            .I(\Lab_UT.scctrl.N_401_0 ));
    Odrv4 I__3010 (
            .O(N__15296),
            .I(\Lab_UT.scctrl.N_401_0 ));
    InMux I__3009 (
            .O(N__15291),
            .I(N__15288));
    LocalMux I__3008 (
            .O(N__15288),
            .I(N__15284));
    InMux I__3007 (
            .O(N__15287),
            .I(N__15281));
    Span4Mux_h I__3006 (
            .O(N__15284),
            .I(N__15278));
    LocalMux I__3005 (
            .O(N__15281),
            .I(N__15275));
    Span4Mux_v I__3004 (
            .O(N__15278),
            .I(N__15272));
    Span4Mux_h I__3003 (
            .O(N__15275),
            .I(N__15269));
    Odrv4 I__3002 (
            .O(N__15272),
            .I(\Lab_UT.scctrl.N_9_0 ));
    Odrv4 I__3001 (
            .O(N__15269),
            .I(\Lab_UT.scctrl.N_9_0 ));
    InMux I__3000 (
            .O(N__15264),
            .I(N__15261));
    LocalMux I__2999 (
            .O(N__15261),
            .I(N__15258));
    Span4Mux_v I__2998 (
            .O(N__15258),
            .I(N__15254));
    InMux I__2997 (
            .O(N__15257),
            .I(N__15251));
    Odrv4 I__2996 (
            .O(N__15254),
            .I(\Lab_UT.scctrl.g0_i_2 ));
    LocalMux I__2995 (
            .O(N__15251),
            .I(\Lab_UT.scctrl.g0_i_2 ));
    CascadeMux I__2994 (
            .O(N__15246),
            .I(\Lab_UT.scctrl.N_170_i_cascade_ ));
    InMux I__2993 (
            .O(N__15243),
            .I(N__15240));
    LocalMux I__2992 (
            .O(N__15240),
            .I(\Lab_UT.scctrl.G_24_i_o6_0_0 ));
    CascadeMux I__2991 (
            .O(N__15237),
            .I(\Lab_UT.scctrl.N_17_i_cascade_ ));
    InMux I__2990 (
            .O(N__15234),
            .I(N__15231));
    LocalMux I__2989 (
            .O(N__15231),
            .I(\Lab_UT.scctrl.N_418_1 ));
    CascadeMux I__2988 (
            .O(N__15228),
            .I(\Lab_UT.scctrl.g0_8_0_cascade_ ));
    InMux I__2987 (
            .O(N__15225),
            .I(N__15222));
    LocalMux I__2986 (
            .O(N__15222),
            .I(\Lab_UT.scctrl.g0_8_2 ));
    CascadeMux I__2985 (
            .O(N__15219),
            .I(N__15215));
    InMux I__2984 (
            .O(N__15218),
            .I(N__15210));
    InMux I__2983 (
            .O(N__15215),
            .I(N__15210));
    LocalMux I__2982 (
            .O(N__15210),
            .I(N__15207));
    Span4Mux_v I__2981 (
            .O(N__15207),
            .I(N__15204));
    Odrv4 I__2980 (
            .O(N__15204),
            .I(\Lab_UT.scctrl.N_444_1 ));
    CascadeMux I__2979 (
            .O(N__15201),
            .I(N__15198));
    InMux I__2978 (
            .O(N__15198),
            .I(N__15190));
    InMux I__2977 (
            .O(N__15197),
            .I(N__15190));
    InMux I__2976 (
            .O(N__15196),
            .I(N__15187));
    InMux I__2975 (
            .O(N__15195),
            .I(N__15184));
    LocalMux I__2974 (
            .O(N__15190),
            .I(N__15177));
    LocalMux I__2973 (
            .O(N__15187),
            .I(N__15172));
    LocalMux I__2972 (
            .O(N__15184),
            .I(N__15172));
    InMux I__2971 (
            .O(N__15183),
            .I(N__15165));
    InMux I__2970 (
            .O(N__15182),
            .I(N__15162));
    InMux I__2969 (
            .O(N__15181),
            .I(N__15159));
    InMux I__2968 (
            .O(N__15180),
            .I(N__15156));
    Span4Mux_v I__2967 (
            .O(N__15177),
            .I(N__15151));
    Span4Mux_v I__2966 (
            .O(N__15172),
            .I(N__15151));
    InMux I__2965 (
            .O(N__15171),
            .I(N__15142));
    InMux I__2964 (
            .O(N__15170),
            .I(N__15142));
    InMux I__2963 (
            .O(N__15169),
            .I(N__15142));
    InMux I__2962 (
            .O(N__15168),
            .I(N__15142));
    LocalMux I__2961 (
            .O(N__15165),
            .I(bu_rx_data_i_1_6));
    LocalMux I__2960 (
            .O(N__15162),
            .I(bu_rx_data_i_1_6));
    LocalMux I__2959 (
            .O(N__15159),
            .I(bu_rx_data_i_1_6));
    LocalMux I__2958 (
            .O(N__15156),
            .I(bu_rx_data_i_1_6));
    Odrv4 I__2957 (
            .O(N__15151),
            .I(bu_rx_data_i_1_6));
    LocalMux I__2956 (
            .O(N__15142),
            .I(bu_rx_data_i_1_6));
    InMux I__2955 (
            .O(N__15129),
            .I(N__15121));
    InMux I__2954 (
            .O(N__15128),
            .I(N__15117));
    InMux I__2953 (
            .O(N__15127),
            .I(N__15113));
    InMux I__2952 (
            .O(N__15126),
            .I(N__15108));
    InMux I__2951 (
            .O(N__15125),
            .I(N__15108));
    InMux I__2950 (
            .O(N__15124),
            .I(N__15101));
    LocalMux I__2949 (
            .O(N__15121),
            .I(N__15098));
    CascadeMux I__2948 (
            .O(N__15120),
            .I(N__15093));
    LocalMux I__2947 (
            .O(N__15117),
            .I(N__15088));
    InMux I__2946 (
            .O(N__15116),
            .I(N__15085));
    LocalMux I__2945 (
            .O(N__15113),
            .I(N__15080));
    LocalMux I__2944 (
            .O(N__15108),
            .I(N__15076));
    InMux I__2943 (
            .O(N__15107),
            .I(N__15064));
    InMux I__2942 (
            .O(N__15106),
            .I(N__15064));
    InMux I__2941 (
            .O(N__15105),
            .I(N__15061));
    InMux I__2940 (
            .O(N__15104),
            .I(N__15058));
    LocalMux I__2939 (
            .O(N__15101),
            .I(N__15053));
    Span4Mux_h I__2938 (
            .O(N__15098),
            .I(N__15053));
    InMux I__2937 (
            .O(N__15097),
            .I(N__15042));
    InMux I__2936 (
            .O(N__15096),
            .I(N__15042));
    InMux I__2935 (
            .O(N__15093),
            .I(N__15042));
    InMux I__2934 (
            .O(N__15092),
            .I(N__15042));
    InMux I__2933 (
            .O(N__15091),
            .I(N__15042));
    Span12Mux_s5_h I__2932 (
            .O(N__15088),
            .I(N__15039));
    LocalMux I__2931 (
            .O(N__15085),
            .I(N__15036));
    InMux I__2930 (
            .O(N__15084),
            .I(N__15033));
    InMux I__2929 (
            .O(N__15083),
            .I(N__15030));
    Span4Mux_v I__2928 (
            .O(N__15080),
            .I(N__15027));
    InMux I__2927 (
            .O(N__15079),
            .I(N__15024));
    Span4Mux_v I__2926 (
            .O(N__15076),
            .I(N__15021));
    InMux I__2925 (
            .O(N__15075),
            .I(N__15018));
    InMux I__2924 (
            .O(N__15074),
            .I(N__15009));
    InMux I__2923 (
            .O(N__15073),
            .I(N__15009));
    InMux I__2922 (
            .O(N__15072),
            .I(N__15009));
    InMux I__2921 (
            .O(N__15071),
            .I(N__15009));
    InMux I__2920 (
            .O(N__15070),
            .I(N__15004));
    InMux I__2919 (
            .O(N__15069),
            .I(N__15004));
    LocalMux I__2918 (
            .O(N__15064),
            .I(N__14999));
    LocalMux I__2917 (
            .O(N__15061),
            .I(N__14999));
    LocalMux I__2916 (
            .O(N__15058),
            .I(N__14994));
    Span4Mux_v I__2915 (
            .O(N__15053),
            .I(N__14994));
    LocalMux I__2914 (
            .O(N__15042),
            .I(N__14991));
    Odrv12 I__2913 (
            .O(N__15039),
            .I(bu_rx_data_4));
    Odrv4 I__2912 (
            .O(N__15036),
            .I(bu_rx_data_4));
    LocalMux I__2911 (
            .O(N__15033),
            .I(bu_rx_data_4));
    LocalMux I__2910 (
            .O(N__15030),
            .I(bu_rx_data_4));
    Odrv4 I__2909 (
            .O(N__15027),
            .I(bu_rx_data_4));
    LocalMux I__2908 (
            .O(N__15024),
            .I(bu_rx_data_4));
    Odrv4 I__2907 (
            .O(N__15021),
            .I(bu_rx_data_4));
    LocalMux I__2906 (
            .O(N__15018),
            .I(bu_rx_data_4));
    LocalMux I__2905 (
            .O(N__15009),
            .I(bu_rx_data_4));
    LocalMux I__2904 (
            .O(N__15004),
            .I(bu_rx_data_4));
    Odrv4 I__2903 (
            .O(N__14999),
            .I(bu_rx_data_4));
    Odrv4 I__2902 (
            .O(N__14994),
            .I(bu_rx_data_4));
    Odrv4 I__2901 (
            .O(N__14991),
            .I(bu_rx_data_4));
    CascadeMux I__2900 (
            .O(N__14964),
            .I(\Lab_UT.scctrl.G_24_i_a6_2_2_cascade_ ));
    InMux I__2899 (
            .O(N__14961),
            .I(N__14958));
    LocalMux I__2898 (
            .O(N__14958),
            .I(N__14955));
    Span4Mux_v I__2897 (
            .O(N__14955),
            .I(N__14952));
    Odrv4 I__2896 (
            .O(N__14952),
            .I(\Lab_UT.scctrl.N_12_3 ));
    CascadeMux I__2895 (
            .O(N__14949),
            .I(N__14945));
    CascadeMux I__2894 (
            .O(N__14948),
            .I(N__14942));
    InMux I__2893 (
            .O(N__14945),
            .I(N__14932));
    InMux I__2892 (
            .O(N__14942),
            .I(N__14927));
    InMux I__2891 (
            .O(N__14941),
            .I(N__14927));
    InMux I__2890 (
            .O(N__14940),
            .I(N__14923));
    CascadeMux I__2889 (
            .O(N__14939),
            .I(N__14920));
    InMux I__2888 (
            .O(N__14938),
            .I(N__14913));
    InMux I__2887 (
            .O(N__14937),
            .I(N__14913));
    InMux I__2886 (
            .O(N__14936),
            .I(N__14913));
    InMux I__2885 (
            .O(N__14935),
            .I(N__14910));
    LocalMux I__2884 (
            .O(N__14932),
            .I(N__14904));
    LocalMux I__2883 (
            .O(N__14927),
            .I(N__14904));
    InMux I__2882 (
            .O(N__14926),
            .I(N__14901));
    LocalMux I__2881 (
            .O(N__14923),
            .I(N__14897));
    InMux I__2880 (
            .O(N__14920),
            .I(N__14894));
    LocalMux I__2879 (
            .O(N__14913),
            .I(N__14891));
    LocalMux I__2878 (
            .O(N__14910),
            .I(N__14888));
    InMux I__2877 (
            .O(N__14909),
            .I(N__14885));
    Span4Mux_h I__2876 (
            .O(N__14904),
            .I(N__14882));
    LocalMux I__2875 (
            .O(N__14901),
            .I(N__14879));
    InMux I__2874 (
            .O(N__14900),
            .I(N__14876));
    Span12Mux_s11_v I__2873 (
            .O(N__14897),
            .I(N__14871));
    LocalMux I__2872 (
            .O(N__14894),
            .I(N__14871));
    Span4Mux_h I__2871 (
            .O(N__14891),
            .I(N__14860));
    Span4Mux_h I__2870 (
            .O(N__14888),
            .I(N__14860));
    LocalMux I__2869 (
            .O(N__14885),
            .I(N__14860));
    Span4Mux_v I__2868 (
            .O(N__14882),
            .I(N__14860));
    Span4Mux_h I__2867 (
            .O(N__14879),
            .I(N__14860));
    LocalMux I__2866 (
            .O(N__14876),
            .I(bu_rx_data_6));
    Odrv12 I__2865 (
            .O(N__14871),
            .I(bu_rx_data_6));
    Odrv4 I__2864 (
            .O(N__14860),
            .I(bu_rx_data_6));
    InMux I__2863 (
            .O(N__14853),
            .I(N__14843));
    InMux I__2862 (
            .O(N__14852),
            .I(N__14843));
    InMux I__2861 (
            .O(N__14851),
            .I(N__14843));
    InMux I__2860 (
            .O(N__14850),
            .I(N__14840));
    LocalMux I__2859 (
            .O(N__14843),
            .I(N__14837));
    LocalMux I__2858 (
            .O(N__14840),
            .I(N__14833));
    Span12Mux_s9_v I__2857 (
            .O(N__14837),
            .I(N__14830));
    InMux I__2856 (
            .O(N__14836),
            .I(N__14827));
    Odrv4 I__2855 (
            .O(N__14833),
            .I(\Lab_UT.scctrl.N_241_i_0 ));
    Odrv12 I__2854 (
            .O(N__14830),
            .I(\Lab_UT.scctrl.N_241_i_0 ));
    LocalMux I__2853 (
            .O(N__14827),
            .I(\Lab_UT.scctrl.N_241_i_0 ));
    InMux I__2852 (
            .O(N__14820),
            .I(N__14817));
    LocalMux I__2851 (
            .O(N__14817),
            .I(\Lab_UT.scctrl.G_24_i_2_0 ));
    InMux I__2850 (
            .O(N__14814),
            .I(N__14811));
    LocalMux I__2849 (
            .O(N__14811),
            .I(\Lab_UT.scctrl.G_24_i_a6_0_2 ));
    CascadeMux I__2848 (
            .O(N__14808),
            .I(\Lab_UT.scctrl.N_5_2_cascade_ ));
    InMux I__2847 (
            .O(N__14805),
            .I(N__14802));
    LocalMux I__2846 (
            .O(N__14802),
            .I(N__14799));
    Odrv12 I__2845 (
            .O(N__14799),
            .I(\Lab_UT.scctrl.next_state_rst_2_1 ));
    InMux I__2844 (
            .O(N__14796),
            .I(N__14793));
    LocalMux I__2843 (
            .O(N__14793),
            .I(\Lab_UT.scctrl.next_state_rst_4_1 ));
    InMux I__2842 (
            .O(N__14790),
            .I(N__14786));
    InMux I__2841 (
            .O(N__14789),
            .I(N__14783));
    LocalMux I__2840 (
            .O(N__14786),
            .I(\Lab_UT.scctrl.G_15_0_a10_1_2 ));
    LocalMux I__2839 (
            .O(N__14783),
            .I(\Lab_UT.scctrl.G_15_0_a10_1_2 ));
    InMux I__2838 (
            .O(N__14778),
            .I(N__14775));
    LocalMux I__2837 (
            .O(N__14775),
            .I(\Lab_UT.scctrl.N_7 ));
    InMux I__2836 (
            .O(N__14772),
            .I(N__14769));
    LocalMux I__2835 (
            .O(N__14769),
            .I(\Lab_UT.scctrl.g0_8_0_0 ));
    InMux I__2834 (
            .O(N__14766),
            .I(N__14763));
    LocalMux I__2833 (
            .O(N__14763),
            .I(N__14759));
    InMux I__2832 (
            .O(N__14762),
            .I(N__14756));
    Span4Mux_v I__2831 (
            .O(N__14759),
            .I(N__14753));
    LocalMux I__2830 (
            .O(N__14756),
            .I(N__14750));
    Odrv4 I__2829 (
            .O(N__14753),
            .I(\Lab_UT.scctrl.N_223_0_0 ));
    Odrv4 I__2828 (
            .O(N__14750),
            .I(\Lab_UT.scctrl.N_223_0_0 ));
    CascadeMux I__2827 (
            .O(N__14745),
            .I(\Lab_UT.scctrl.N_419_0_cascade_ ));
    InMux I__2826 (
            .O(N__14742),
            .I(N__14739));
    LocalMux I__2825 (
            .O(N__14739),
            .I(N__14736));
    Span4Mux_h I__2824 (
            .O(N__14736),
            .I(N__14733));
    Odrv4 I__2823 (
            .O(N__14733),
            .I(\Lab_UT.scctrl.g1 ));
    CascadeMux I__2822 (
            .O(N__14730),
            .I(N__14727));
    InMux I__2821 (
            .O(N__14727),
            .I(N__14724));
    LocalMux I__2820 (
            .O(N__14724),
            .I(N__14721));
    Span4Mux_v I__2819 (
            .O(N__14721),
            .I(N__14718));
    Odrv4 I__2818 (
            .O(N__14718),
            .I(\Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_0_3 ));
    CascadeMux I__2817 (
            .O(N__14715),
            .I(\Lab_UT.scctrl.g0_2_0_0_a3_2_cascade_ ));
    InMux I__2816 (
            .O(N__14712),
            .I(N__14709));
    LocalMux I__2815 (
            .O(N__14709),
            .I(N__14706));
    Odrv12 I__2814 (
            .O(N__14706),
            .I(\Lab_UT.scctrl.G_24_i_a3_3 ));
    CascadeMux I__2813 (
            .O(N__14703),
            .I(\Lab_UT.scctrl.G_24_i_a3_5_cascade_ ));
    InMux I__2812 (
            .O(N__14700),
            .I(N__14697));
    LocalMux I__2811 (
            .O(N__14697),
            .I(\Lab_UT.scctrl.G_24_i_a3_0_3 ));
    CascadeMux I__2810 (
            .O(N__14694),
            .I(N__14691));
    InMux I__2809 (
            .O(N__14691),
            .I(N__14688));
    LocalMux I__2808 (
            .O(N__14688),
            .I(\Lab_UT.scctrl.G_24_i_a3_0_1 ));
    InMux I__2807 (
            .O(N__14685),
            .I(N__14682));
    LocalMux I__2806 (
            .O(N__14682),
            .I(N__14679));
    Odrv4 I__2805 (
            .O(N__14679),
            .I(\Lab_UT.scctrl.N_15 ));
    CascadeMux I__2804 (
            .O(N__14676),
            .I(N__14673));
    InMux I__2803 (
            .O(N__14673),
            .I(N__14670));
    LocalMux I__2802 (
            .O(N__14670),
            .I(\Lab_UT.scctrl.next_state_rst_0_3_tz_0 ));
    CascadeMux I__2801 (
            .O(N__14667),
            .I(\Lab_UT.scctrl.g0_0_4_cascade_ ));
    CascadeMux I__2800 (
            .O(N__14664),
            .I(\Lab_UT.scctrl.next_state_rst_cascade_ ));
    CascadeMux I__2799 (
            .O(N__14661),
            .I(N__14657));
    CascadeMux I__2798 (
            .O(N__14660),
            .I(N__14654));
    InMux I__2797 (
            .O(N__14657),
            .I(N__14647));
    InMux I__2796 (
            .O(N__14654),
            .I(N__14647));
    InMux I__2795 (
            .O(N__14653),
            .I(N__14644));
    InMux I__2794 (
            .O(N__14652),
            .I(N__14641));
    LocalMux I__2793 (
            .O(N__14647),
            .I(N__14638));
    LocalMux I__2792 (
            .O(N__14644),
            .I(N__14623));
    LocalMux I__2791 (
            .O(N__14641),
            .I(N__14623));
    Span4Mux_h I__2790 (
            .O(N__14638),
            .I(N__14623));
    InMux I__2789 (
            .O(N__14637),
            .I(N__14612));
    InMux I__2788 (
            .O(N__14636),
            .I(N__14612));
    InMux I__2787 (
            .O(N__14635),
            .I(N__14612));
    InMux I__2786 (
            .O(N__14634),
            .I(N__14612));
    InMux I__2785 (
            .O(N__14633),
            .I(N__14612));
    InMux I__2784 (
            .O(N__14632),
            .I(N__14609));
    InMux I__2783 (
            .O(N__14631),
            .I(N__14604));
    InMux I__2782 (
            .O(N__14630),
            .I(N__14604));
    Span4Mux_v I__2781 (
            .O(N__14623),
            .I(N__14599));
    LocalMux I__2780 (
            .O(N__14612),
            .I(N__14599));
    LocalMux I__2779 (
            .O(N__14609),
            .I(N__14596));
    LocalMux I__2778 (
            .O(N__14604),
            .I(N__14593));
    Span4Mux_v I__2777 (
            .O(N__14599),
            .I(N__14589));
    Span4Mux_h I__2776 (
            .O(N__14596),
            .I(N__14584));
    Span4Mux_v I__2775 (
            .O(N__14593),
            .I(N__14584));
    InMux I__2774 (
            .O(N__14592),
            .I(N__14581));
    Odrv4 I__2773 (
            .O(N__14589),
            .I(\Lab_UT.scctrl.state_i_1_0_rep2 ));
    Odrv4 I__2772 (
            .O(N__14584),
            .I(\Lab_UT.scctrl.state_i_1_0_rep2 ));
    LocalMux I__2771 (
            .O(N__14581),
            .I(\Lab_UT.scctrl.state_i_1_0_rep2 ));
    CascadeMux I__2770 (
            .O(N__14574),
            .I(\Lab_UT.scctrl.N_299_i_0_cascade_ ));
    InMux I__2769 (
            .O(N__14571),
            .I(N__14567));
    InMux I__2768 (
            .O(N__14570),
            .I(N__14564));
    LocalMux I__2767 (
            .O(N__14567),
            .I(N__14559));
    LocalMux I__2766 (
            .O(N__14564),
            .I(N__14559));
    Odrv4 I__2765 (
            .O(N__14559),
            .I(\Lab_UT.scctrl.N_4 ));
    InMux I__2764 (
            .O(N__14556),
            .I(N__14553));
    LocalMux I__2763 (
            .O(N__14553),
            .I(\Lab_UT.scctrl.N_240_reti ));
    InMux I__2762 (
            .O(N__14550),
            .I(N__14547));
    LocalMux I__2761 (
            .O(N__14547),
            .I(\Lab_UT.scctrl.N_419_1 ));
    CascadeMux I__2760 (
            .O(N__14544),
            .I(\Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_2_3_cascade_ ));
    CascadeMux I__2759 (
            .O(N__14541),
            .I(N__14538));
    InMux I__2758 (
            .O(N__14538),
            .I(N__14535));
    LocalMux I__2757 (
            .O(N__14535),
            .I(N__14532));
    Odrv4 I__2756 (
            .O(N__14532),
            .I(\Lab_UT.scctrl.g0_0_0 ));
    InMux I__2755 (
            .O(N__14529),
            .I(N__14523));
    InMux I__2754 (
            .O(N__14528),
            .I(N__14511));
    InMux I__2753 (
            .O(N__14527),
            .I(N__14507));
    InMux I__2752 (
            .O(N__14526),
            .I(N__14504));
    LocalMux I__2751 (
            .O(N__14523),
            .I(N__14501));
    InMux I__2750 (
            .O(N__14522),
            .I(N__14498));
    InMux I__2749 (
            .O(N__14521),
            .I(N__14493));
    InMux I__2748 (
            .O(N__14520),
            .I(N__14493));
    InMux I__2747 (
            .O(N__14519),
            .I(N__14486));
    InMux I__2746 (
            .O(N__14518),
            .I(N__14486));
    InMux I__2745 (
            .O(N__14517),
            .I(N__14486));
    InMux I__2744 (
            .O(N__14516),
            .I(N__14483));
    InMux I__2743 (
            .O(N__14515),
            .I(N__14479));
    InMux I__2742 (
            .O(N__14514),
            .I(N__14476));
    LocalMux I__2741 (
            .O(N__14511),
            .I(N__14471));
    InMux I__2740 (
            .O(N__14510),
            .I(N__14465));
    LocalMux I__2739 (
            .O(N__14507),
            .I(N__14460));
    LocalMux I__2738 (
            .O(N__14504),
            .I(N__14460));
    Span4Mux_v I__2737 (
            .O(N__14501),
            .I(N__14455));
    LocalMux I__2736 (
            .O(N__14498),
            .I(N__14455));
    LocalMux I__2735 (
            .O(N__14493),
            .I(N__14450));
    LocalMux I__2734 (
            .O(N__14486),
            .I(N__14450));
    LocalMux I__2733 (
            .O(N__14483),
            .I(N__14447));
    InMux I__2732 (
            .O(N__14482),
            .I(N__14444));
    LocalMux I__2731 (
            .O(N__14479),
            .I(N__14441));
    LocalMux I__2730 (
            .O(N__14476),
            .I(N__14438));
    InMux I__2729 (
            .O(N__14475),
            .I(N__14433));
    InMux I__2728 (
            .O(N__14474),
            .I(N__14433));
    Span4Mux_h I__2727 (
            .O(N__14471),
            .I(N__14430));
    InMux I__2726 (
            .O(N__14470),
            .I(N__14425));
    InMux I__2725 (
            .O(N__14469),
            .I(N__14425));
    InMux I__2724 (
            .O(N__14468),
            .I(N__14422));
    LocalMux I__2723 (
            .O(N__14465),
            .I(N__14419));
    Span4Mux_v I__2722 (
            .O(N__14460),
            .I(N__14412));
    Span4Mux_h I__2721 (
            .O(N__14455),
            .I(N__14412));
    Span4Mux_h I__2720 (
            .O(N__14450),
            .I(N__14412));
    Span4Mux_h I__2719 (
            .O(N__14447),
            .I(N__14407));
    LocalMux I__2718 (
            .O(N__14444),
            .I(N__14407));
    Span4Mux_h I__2717 (
            .O(N__14441),
            .I(N__14400));
    Span4Mux_v I__2716 (
            .O(N__14438),
            .I(N__14400));
    LocalMux I__2715 (
            .O(N__14433),
            .I(N__14400));
    Odrv4 I__2714 (
            .O(N__14430),
            .I(bu_rx_data_7));
    LocalMux I__2713 (
            .O(N__14425),
            .I(bu_rx_data_7));
    LocalMux I__2712 (
            .O(N__14422),
            .I(bu_rx_data_7));
    Odrv12 I__2711 (
            .O(N__14419),
            .I(bu_rx_data_7));
    Odrv4 I__2710 (
            .O(N__14412),
            .I(bu_rx_data_7));
    Odrv4 I__2709 (
            .O(N__14407),
            .I(bu_rx_data_7));
    Odrv4 I__2708 (
            .O(N__14400),
            .I(bu_rx_data_7));
    InMux I__2707 (
            .O(N__14385),
            .I(N__14375));
    InMux I__2706 (
            .O(N__14384),
            .I(N__14375));
    InMux I__2705 (
            .O(N__14383),
            .I(N__14367));
    InMux I__2704 (
            .O(N__14382),
            .I(N__14361));
    InMux I__2703 (
            .O(N__14381),
            .I(N__14361));
    InMux I__2702 (
            .O(N__14380),
            .I(N__14358));
    LocalMux I__2701 (
            .O(N__14375),
            .I(N__14355));
    InMux I__2700 (
            .O(N__14374),
            .I(N__14348));
    InMux I__2699 (
            .O(N__14373),
            .I(N__14348));
    InMux I__2698 (
            .O(N__14372),
            .I(N__14348));
    InMux I__2697 (
            .O(N__14371),
            .I(N__14345));
    InMux I__2696 (
            .O(N__14370),
            .I(N__14342));
    LocalMux I__2695 (
            .O(N__14367),
            .I(N__14339));
    InMux I__2694 (
            .O(N__14366),
            .I(N__14335));
    LocalMux I__2693 (
            .O(N__14361),
            .I(N__14332));
    LocalMux I__2692 (
            .O(N__14358),
            .I(N__14323));
    Span4Mux_v I__2691 (
            .O(N__14355),
            .I(N__14323));
    LocalMux I__2690 (
            .O(N__14348),
            .I(N__14323));
    LocalMux I__2689 (
            .O(N__14345),
            .I(N__14323));
    LocalMux I__2688 (
            .O(N__14342),
            .I(N__14320));
    Span4Mux_v I__2687 (
            .O(N__14339),
            .I(N__14317));
    InMux I__2686 (
            .O(N__14338),
            .I(N__14314));
    LocalMux I__2685 (
            .O(N__14335),
            .I(N__14311));
    Span4Mux_v I__2684 (
            .O(N__14332),
            .I(N__14306));
    Span4Mux_h I__2683 (
            .O(N__14323),
            .I(N__14306));
    Span4Mux_h I__2682 (
            .O(N__14320),
            .I(N__14299));
    Span4Mux_h I__2681 (
            .O(N__14317),
            .I(N__14299));
    LocalMux I__2680 (
            .O(N__14314),
            .I(N__14299));
    Odrv4 I__2679 (
            .O(N__14311),
            .I(N_232));
    Odrv4 I__2678 (
            .O(N__14306),
            .I(N_232));
    Odrv4 I__2677 (
            .O(N__14299),
            .I(N_232));
    InMux I__2676 (
            .O(N__14292),
            .I(N__14289));
    LocalMux I__2675 (
            .O(N__14289),
            .I(N__14286));
    Span4Mux_v I__2674 (
            .O(N__14286),
            .I(N__14283));
    Odrv4 I__2673 (
            .O(N__14283),
            .I(\Lab_UT.scctrl.g0_2_0 ));
    CascadeMux I__2672 (
            .O(N__14280),
            .I(\Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_1_3_cascade_ ));
    InMux I__2671 (
            .O(N__14277),
            .I(N__14274));
    LocalMux I__2670 (
            .O(N__14274),
            .I(N__14271));
    Odrv12 I__2669 (
            .O(N__14271),
            .I(\Lab_UT.scctrl.next_state_0_0 ));
    InMux I__2668 (
            .O(N__14268),
            .I(N__14265));
    LocalMux I__2667 (
            .O(N__14265),
            .I(\Lab_UT.scctrl.g0_1_i_0 ));
    CascadeMux I__2666 (
            .O(N__14262),
            .I(\Lab_UT.scctrl.g0_1_i_2_cascade_ ));
    InMux I__2665 (
            .O(N__14259),
            .I(N__14256));
    LocalMux I__2664 (
            .O(N__14256),
            .I(\Lab_UT.scctrl.g0_1_i_4 ));
    InMux I__2663 (
            .O(N__14253),
            .I(N__14250));
    LocalMux I__2662 (
            .O(N__14250),
            .I(N__14247));
    Odrv4 I__2661 (
            .O(N__14247),
            .I(\Lab_UT.scctrl.next_state_rst_2_0 ));
    CascadeMux I__2660 (
            .O(N__14244),
            .I(\Lab_UT.scctrl.G_24_i_a3_0_cascade_ ));
    InMux I__2659 (
            .O(N__14241),
            .I(N__14238));
    LocalMux I__2658 (
            .O(N__14238),
            .I(\Lab_UT.scctrl.N_8 ));
    CascadeMux I__2657 (
            .O(N__14235),
            .I(\Lab_UT.scctrl.N_290_2_cascade_ ));
    InMux I__2656 (
            .O(N__14232),
            .I(N__14229));
    LocalMux I__2655 (
            .O(N__14229),
            .I(\Lab_UT.scctrl.N_8_3 ));
    InMux I__2654 (
            .O(N__14226),
            .I(N__14223));
    LocalMux I__2653 (
            .O(N__14223),
            .I(\Lab_UT.scctrl.g0_1_2_0 ));
    CascadeMux I__2652 (
            .O(N__14220),
            .I(\Lab_UT.scctrl.g3_cascade_ ));
    InMux I__2651 (
            .O(N__14217),
            .I(N__14214));
    LocalMux I__2650 (
            .O(N__14214),
            .I(\Lab_UT.scctrl.g0_1_4 ));
    CascadeMux I__2649 (
            .O(N__14211),
            .I(\Lab_UT.scctrl.next_state_rst_1_cascade_ ));
    InMux I__2648 (
            .O(N__14208),
            .I(N__14205));
    LocalMux I__2647 (
            .O(N__14205),
            .I(N__14202));
    Span4Mux_v I__2646 (
            .O(N__14202),
            .I(N__14199));
    Odrv4 I__2645 (
            .O(N__14199),
            .I(\Lab_UT.scctrl.g0_i_0 ));
    CascadeMux I__2644 (
            .O(N__14196),
            .I(N__14193));
    InMux I__2643 (
            .O(N__14193),
            .I(N__14190));
    LocalMux I__2642 (
            .O(N__14190),
            .I(N__14187));
    Odrv4 I__2641 (
            .O(N__14187),
            .I(\Lab_UT.scctrl.g3_0 ));
    CascadeMux I__2640 (
            .O(N__14184),
            .I(\Lab_UT.scctrl.next_state_rst_0_7_cascade_ ));
    InMux I__2639 (
            .O(N__14181),
            .I(N__14178));
    LocalMux I__2638 (
            .O(N__14178),
            .I(\Lab_UT.scctrl.N_10 ));
    CascadeMux I__2637 (
            .O(N__14175),
            .I(\Lab_UT.scctrl.g1_0_4_cascade_ ));
    InMux I__2636 (
            .O(N__14172),
            .I(N__14169));
    LocalMux I__2635 (
            .O(N__14169),
            .I(\Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_3 ));
    CascadeMux I__2634 (
            .O(N__14166),
            .I(\Lab_UT.scctrl.N_290_cascade_ ));
    CascadeMux I__2633 (
            .O(N__14163),
            .I(\Lab_UT.scctrl.N_9_cascade_ ));
    InMux I__2632 (
            .O(N__14160),
            .I(N__14157));
    LocalMux I__2631 (
            .O(N__14157),
            .I(\Lab_UT.scctrl.g0_9_0 ));
    InMux I__2630 (
            .O(N__14154),
            .I(N__14151));
    LocalMux I__2629 (
            .O(N__14151),
            .I(N__14147));
    CascadeMux I__2628 (
            .O(N__14150),
            .I(N__14144));
    Span12Mux_v I__2627 (
            .O(N__14147),
            .I(N__14141));
    InMux I__2626 (
            .O(N__14144),
            .I(N__14138));
    Odrv12 I__2625 (
            .O(N__14141),
            .I(\Lab_UT.scdp.key1_7 ));
    LocalMux I__2624 (
            .O(N__14138),
            .I(\Lab_UT.scdp.key1_7 ));
    CascadeMux I__2623 (
            .O(N__14133),
            .I(N__14129));
    InMux I__2622 (
            .O(N__14132),
            .I(N__14126));
    InMux I__2621 (
            .O(N__14129),
            .I(N__14123));
    LocalMux I__2620 (
            .O(N__14126),
            .I(\Lab_UT.scdp.key1_0 ));
    LocalMux I__2619 (
            .O(N__14123),
            .I(\Lab_UT.scdp.key1_0 ));
    CascadeMux I__2618 (
            .O(N__14118),
            .I(N__14114));
    InMux I__2617 (
            .O(N__14117),
            .I(N__14111));
    InMux I__2616 (
            .O(N__14114),
            .I(N__14108));
    LocalMux I__2615 (
            .O(N__14111),
            .I(\Lab_UT.scdp.key1_3 ));
    LocalMux I__2614 (
            .O(N__14108),
            .I(\Lab_UT.scdp.key1_3 ));
    InMux I__2613 (
            .O(N__14103),
            .I(N__14100));
    LocalMux I__2612 (
            .O(N__14100),
            .I(N__14096));
    InMux I__2611 (
            .O(N__14099),
            .I(N__14093));
    Odrv4 I__2610 (
            .O(N__14096),
            .I(\Lab_UT.scdp.key2_6 ));
    LocalMux I__2609 (
            .O(N__14093),
            .I(\Lab_UT.scdp.key2_6 ));
    CascadeMux I__2608 (
            .O(N__14088),
            .I(N__14084));
    InMux I__2607 (
            .O(N__14087),
            .I(N__14081));
    InMux I__2606 (
            .O(N__14084),
            .I(N__14078));
    LocalMux I__2605 (
            .O(N__14081),
            .I(\Lab_UT.scdp.key2_4 ));
    LocalMux I__2604 (
            .O(N__14078),
            .I(\Lab_UT.scdp.key2_4 ));
    CascadeMux I__2603 (
            .O(N__14073),
            .I(N__14069));
    InMux I__2602 (
            .O(N__14072),
            .I(N__14066));
    InMux I__2601 (
            .O(N__14069),
            .I(N__14063));
    LocalMux I__2600 (
            .O(N__14066),
            .I(\Lab_UT.scdp.key2_2 ));
    LocalMux I__2599 (
            .O(N__14063),
            .I(\Lab_UT.scdp.key2_2 ));
    InMux I__2598 (
            .O(N__14058),
            .I(N__14055));
    LocalMux I__2597 (
            .O(N__14055),
            .I(N__14052));
    Span4Mux_s2_v I__2596 (
            .O(N__14052),
            .I(N__14048));
    InMux I__2595 (
            .O(N__14051),
            .I(N__14045));
    Odrv4 I__2594 (
            .O(N__14048),
            .I(\Lab_UT.scdp.key1_2 ));
    LocalMux I__2593 (
            .O(N__14045),
            .I(\Lab_UT.scdp.key1_2 ));
    InMux I__2592 (
            .O(N__14040),
            .I(N__14037));
    LocalMux I__2591 (
            .O(N__14037),
            .I(N__14033));
    CascadeMux I__2590 (
            .O(N__14036),
            .I(N__14030));
    Span4Mux_h I__2589 (
            .O(N__14033),
            .I(N__14027));
    InMux I__2588 (
            .O(N__14030),
            .I(N__14024));
    Odrv4 I__2587 (
            .O(N__14027),
            .I(\Lab_UT.scdp.key2_5 ));
    LocalMux I__2586 (
            .O(N__14024),
            .I(\Lab_UT.scdp.key2_5 ));
    CascadeMux I__2585 (
            .O(N__14019),
            .I(N__14015));
    InMux I__2584 (
            .O(N__14018),
            .I(N__14012));
    InMux I__2583 (
            .O(N__14015),
            .I(N__14009));
    LocalMux I__2582 (
            .O(N__14012),
            .I(\Lab_UT.scdp.key1_4 ));
    LocalMux I__2581 (
            .O(N__14009),
            .I(\Lab_UT.scdp.key1_4 ));
    CascadeMux I__2580 (
            .O(N__14004),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_cascade_ ));
    CascadeMux I__2579 (
            .O(N__14001),
            .I(N__13997));
    InMux I__2578 (
            .O(N__14000),
            .I(N__13994));
    InMux I__2577 (
            .O(N__13997),
            .I(N__13991));
    LocalMux I__2576 (
            .O(N__13994),
            .I(N__13988));
    LocalMux I__2575 (
            .O(N__13991),
            .I(N__13985));
    Span4Mux_h I__2574 (
            .O(N__13988),
            .I(N__13981));
    Span4Mux_v I__2573 (
            .O(N__13985),
            .I(N__13978));
    InMux I__2572 (
            .O(N__13984),
            .I(N__13975));
    Odrv4 I__2571 (
            .O(N__13981),
            .I(\Lab_UT.scctrl.N_351 ));
    Odrv4 I__2570 (
            .O(N__13978),
            .I(\Lab_UT.scctrl.N_351 ));
    LocalMux I__2569 (
            .O(N__13975),
            .I(\Lab_UT.scctrl.N_351 ));
    InMux I__2568 (
            .O(N__13968),
            .I(N__13965));
    LocalMux I__2567 (
            .O(N__13965),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0 ));
    CascadeMux I__2566 (
            .O(N__13962),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_0_0_cascade_ ));
    InMux I__2565 (
            .O(N__13959),
            .I(N__13956));
    LocalMux I__2564 (
            .O(N__13956),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_2 ));
    InMux I__2563 (
            .O(N__13953),
            .I(N__13950));
    LocalMux I__2562 (
            .O(N__13950),
            .I(N__13947));
    Odrv12 I__2561 (
            .O(N__13947),
            .I(\Lab_UT.scctrl.N_6_2 ));
    InMux I__2560 (
            .O(N__13944),
            .I(N__13941));
    LocalMux I__2559 (
            .O(N__13941),
            .I(\Lab_UT.scctrl.g0_8_1_0 ));
    InMux I__2558 (
            .O(N__13938),
            .I(N__13935));
    LocalMux I__2557 (
            .O(N__13935),
            .I(N__13932));
    Odrv4 I__2556 (
            .O(N__13932),
            .I(\Lab_UT.scctrl.N_404_2 ));
    CascadeMux I__2555 (
            .O(N__13929),
            .I(\Lab_UT.scctrl.g0_8_1_cascade_ ));
    InMux I__2554 (
            .O(N__13926),
            .I(N__13922));
    CascadeMux I__2553 (
            .O(N__13925),
            .I(N__13919));
    LocalMux I__2552 (
            .O(N__13922),
            .I(N__13916));
    InMux I__2551 (
            .O(N__13919),
            .I(N__13913));
    Odrv12 I__2550 (
            .O(N__13916),
            .I(\Lab_UT.scdp.key1_6 ));
    LocalMux I__2549 (
            .O(N__13913),
            .I(\Lab_UT.scdp.key1_6 ));
    CascadeMux I__2548 (
            .O(N__13908),
            .I(\Lab_UT.N_100_i_cascade_ ));
    CEMux I__2547 (
            .O(N__13905),
            .I(N__13902));
    LocalMux I__2546 (
            .O(N__13902),
            .I(N__13899));
    Odrv12 I__2545 (
            .O(N__13899),
            .I(\Lab_UT.scdp.u2.N_100_i_0 ));
    CascadeMux I__2544 (
            .O(N__13896),
            .I(\Lab_UT.scctrl.N_13_0_cascade_ ));
    CascadeMux I__2543 (
            .O(N__13893),
            .I(\Lab_UT.scctrl.N_404_3_cascade_ ));
    InMux I__2542 (
            .O(N__13890),
            .I(N__13877));
    InMux I__2541 (
            .O(N__13889),
            .I(N__13877));
    InMux I__2540 (
            .O(N__13888),
            .I(N__13877));
    InMux I__2539 (
            .O(N__13887),
            .I(N__13877));
    InMux I__2538 (
            .O(N__13886),
            .I(N__13874));
    LocalMux I__2537 (
            .O(N__13877),
            .I(\buart.Z_rx.N_80 ));
    LocalMux I__2536 (
            .O(N__13874),
            .I(\buart.Z_rx.N_80 ));
    InMux I__2535 (
            .O(N__13869),
            .I(N__13866));
    LocalMux I__2534 (
            .O(N__13866),
            .I(N__13862));
    InMux I__2533 (
            .O(N__13865),
            .I(N__13854));
    Span4Mux_h I__2532 (
            .O(N__13862),
            .I(N__13851));
    InMux I__2531 (
            .O(N__13861),
            .I(N__13848));
    InMux I__2530 (
            .O(N__13860),
            .I(N__13843));
    InMux I__2529 (
            .O(N__13859),
            .I(N__13843));
    InMux I__2528 (
            .O(N__13858),
            .I(N__13838));
    InMux I__2527 (
            .O(N__13857),
            .I(N__13838));
    LocalMux I__2526 (
            .O(N__13854),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    Odrv4 I__2525 (
            .O(N__13851),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    LocalMux I__2524 (
            .O(N__13848),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    LocalMux I__2523 (
            .O(N__13843),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    LocalMux I__2522 (
            .O(N__13838),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    CascadeMux I__2521 (
            .O(N__13827),
            .I(N__13823));
    CascadeMux I__2520 (
            .O(N__13826),
            .I(N__13817));
    InMux I__2519 (
            .O(N__13823),
            .I(N__13814));
    InMux I__2518 (
            .O(N__13822),
            .I(N__13811));
    InMux I__2517 (
            .O(N__13821),
            .I(N__13808));
    InMux I__2516 (
            .O(N__13820),
            .I(N__13803));
    InMux I__2515 (
            .O(N__13817),
            .I(N__13803));
    LocalMux I__2514 (
            .O(N__13814),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__2513 (
            .O(N__13811),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__2512 (
            .O(N__13808),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__2511 (
            .O(N__13803),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    InMux I__2510 (
            .O(N__13794),
            .I(N__13787));
    InMux I__2509 (
            .O(N__13793),
            .I(N__13784));
    InMux I__2508 (
            .O(N__13792),
            .I(N__13781));
    InMux I__2507 (
            .O(N__13791),
            .I(N__13776));
    InMux I__2506 (
            .O(N__13790),
            .I(N__13776));
    LocalMux I__2505 (
            .O(N__13787),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    LocalMux I__2504 (
            .O(N__13784),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    LocalMux I__2503 (
            .O(N__13781),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    LocalMux I__2502 (
            .O(N__13776),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    InMux I__2501 (
            .O(N__13767),
            .I(N__13757));
    InMux I__2500 (
            .O(N__13766),
            .I(N__13757));
    InMux I__2499 (
            .O(N__13765),
            .I(N__13757));
    InMux I__2498 (
            .O(N__13764),
            .I(N__13754));
    LocalMux I__2497 (
            .O(N__13757),
            .I(buart__rx_N_86_i_0_o2_1_0));
    LocalMux I__2496 (
            .O(N__13754),
            .I(buart__rx_N_86_i_0_o2_1_0));
    InMux I__2495 (
            .O(N__13749),
            .I(N__13744));
    InMux I__2494 (
            .O(N__13748),
            .I(N__13739));
    InMux I__2493 (
            .O(N__13747),
            .I(N__13739));
    LocalMux I__2492 (
            .O(N__13744),
            .I(N__13736));
    LocalMux I__2491 (
            .O(N__13739),
            .I(\Lab_UT.N_252 ));
    Odrv4 I__2490 (
            .O(N__13736),
            .I(\Lab_UT.N_252 ));
    CascadeMux I__2489 (
            .O(N__13731),
            .I(N__13727));
    CascadeMux I__2488 (
            .O(N__13730),
            .I(N__13718));
    InMux I__2487 (
            .O(N__13727),
            .I(N__13713));
    InMux I__2486 (
            .O(N__13726),
            .I(N__13710));
    InMux I__2485 (
            .O(N__13725),
            .I(N__13703));
    InMux I__2484 (
            .O(N__13724),
            .I(N__13703));
    InMux I__2483 (
            .O(N__13723),
            .I(N__13703));
    InMux I__2482 (
            .O(N__13722),
            .I(N__13694));
    InMux I__2481 (
            .O(N__13721),
            .I(N__13694));
    InMux I__2480 (
            .O(N__13718),
            .I(N__13694));
    InMux I__2479 (
            .O(N__13717),
            .I(N__13694));
    InMux I__2478 (
            .O(N__13716),
            .I(N__13691));
    LocalMux I__2477 (
            .O(N__13713),
            .I(buart__rx_bitcount_4));
    LocalMux I__2476 (
            .O(N__13710),
            .I(buart__rx_bitcount_4));
    LocalMux I__2475 (
            .O(N__13703),
            .I(buart__rx_bitcount_4));
    LocalMux I__2474 (
            .O(N__13694),
            .I(buart__rx_bitcount_4));
    LocalMux I__2473 (
            .O(N__13691),
            .I(buart__rx_bitcount_4));
    CascadeMux I__2472 (
            .O(N__13680),
            .I(buart__rx_N_86_i_0_o2_1_0_cascade_));
    InMux I__2471 (
            .O(N__13677),
            .I(N__13664));
    InMux I__2470 (
            .O(N__13676),
            .I(N__13661));
    InMux I__2469 (
            .O(N__13675),
            .I(N__13658));
    InMux I__2468 (
            .O(N__13674),
            .I(N__13649));
    InMux I__2467 (
            .O(N__13673),
            .I(N__13649));
    InMux I__2466 (
            .O(N__13672),
            .I(N__13649));
    InMux I__2465 (
            .O(N__13671),
            .I(N__13649));
    InMux I__2464 (
            .O(N__13670),
            .I(N__13646));
    InMux I__2463 (
            .O(N__13669),
            .I(N__13639));
    InMux I__2462 (
            .O(N__13668),
            .I(N__13639));
    InMux I__2461 (
            .O(N__13667),
            .I(N__13639));
    LocalMux I__2460 (
            .O(N__13664),
            .I(buart__rx_bitcount_1));
    LocalMux I__2459 (
            .O(N__13661),
            .I(buart__rx_bitcount_1));
    LocalMux I__2458 (
            .O(N__13658),
            .I(buart__rx_bitcount_1));
    LocalMux I__2457 (
            .O(N__13649),
            .I(buart__rx_bitcount_1));
    LocalMux I__2456 (
            .O(N__13646),
            .I(buart__rx_bitcount_1));
    LocalMux I__2455 (
            .O(N__13639),
            .I(buart__rx_bitcount_1));
    InMux I__2454 (
            .O(N__13626),
            .I(N__13623));
    LocalMux I__2453 (
            .O(N__13623),
            .I(N__13620));
    Span4Mux_h I__2452 (
            .O(N__13620),
            .I(N__13617));
    Odrv4 I__2451 (
            .O(N__13617),
            .I(\Lab_UT.scctrl.r4.delay4 ));
    InMux I__2450 (
            .O(N__13614),
            .I(N__13611));
    LocalMux I__2449 (
            .O(N__13611),
            .I(N__13607));
    InMux I__2448 (
            .O(N__13610),
            .I(N__13604));
    Span4Mux_h I__2447 (
            .O(N__13607),
            .I(N__13601));
    LocalMux I__2446 (
            .O(N__13604),
            .I(\Lab_UT.scctrl.delay3 ));
    Odrv4 I__2445 (
            .O(N__13601),
            .I(\Lab_UT.scctrl.delay3 ));
    InMux I__2444 (
            .O(N__13596),
            .I(N__13593));
    LocalMux I__2443 (
            .O(N__13593),
            .I(\Lab_UT.scctrl.delay1 ));
    InMux I__2442 (
            .O(N__13590),
            .I(N__13587));
    LocalMux I__2441 (
            .O(N__13587),
            .I(\Lab_UT.scctrl.delay2 ));
    InMux I__2440 (
            .O(N__13584),
            .I(N__13581));
    LocalMux I__2439 (
            .O(N__13581),
            .I(\Lab_UT.scctrl.N_384 ));
    InMux I__2438 (
            .O(N__13578),
            .I(N__13572));
    InMux I__2437 (
            .O(N__13577),
            .I(N__13572));
    LocalMux I__2436 (
            .O(N__13572),
            .I(N__13569));
    Odrv12 I__2435 (
            .O(N__13569),
            .I(\Lab_UT.scctrl.N_385 ));
    CascadeMux I__2434 (
            .O(N__13566),
            .I(\Lab_UT.scctrl.N_384_cascade_ ));
    InMux I__2433 (
            .O(N__13563),
            .I(N__13559));
    InMux I__2432 (
            .O(N__13562),
            .I(N__13556));
    LocalMux I__2431 (
            .O(N__13559),
            .I(buart__rx_shifter_0_fast_2));
    LocalMux I__2430 (
            .O(N__13556),
            .I(buart__rx_shifter_0_fast_2));
    InMux I__2429 (
            .O(N__13551),
            .I(N__13542));
    CascadeMux I__2428 (
            .O(N__13550),
            .I(N__13538));
    CascadeMux I__2427 (
            .O(N__13549),
            .I(N__13534));
    InMux I__2426 (
            .O(N__13548),
            .I(N__13531));
    InMux I__2425 (
            .O(N__13547),
            .I(N__13524));
    InMux I__2424 (
            .O(N__13546),
            .I(N__13524));
    InMux I__2423 (
            .O(N__13545),
            .I(N__13524));
    LocalMux I__2422 (
            .O(N__13542),
            .I(N__13521));
    InMux I__2421 (
            .O(N__13541),
            .I(N__13518));
    InMux I__2420 (
            .O(N__13538),
            .I(N__13510));
    InMux I__2419 (
            .O(N__13537),
            .I(N__13510));
    InMux I__2418 (
            .O(N__13534),
            .I(N__13510));
    LocalMux I__2417 (
            .O(N__13531),
            .I(N__13505));
    LocalMux I__2416 (
            .O(N__13524),
            .I(N__13502));
    Span4Mux_v I__2415 (
            .O(N__13521),
            .I(N__13498));
    LocalMux I__2414 (
            .O(N__13518),
            .I(N__13495));
    CascadeMux I__2413 (
            .O(N__13517),
            .I(N__13491));
    LocalMux I__2412 (
            .O(N__13510),
            .I(N__13488));
    InMux I__2411 (
            .O(N__13509),
            .I(N__13483));
    InMux I__2410 (
            .O(N__13508),
            .I(N__13483));
    Span4Mux_v I__2409 (
            .O(N__13505),
            .I(N__13478));
    Span4Mux_v I__2408 (
            .O(N__13502),
            .I(N__13478));
    InMux I__2407 (
            .O(N__13501),
            .I(N__13475));
    Span4Mux_h I__2406 (
            .O(N__13498),
            .I(N__13470));
    Span4Mux_v I__2405 (
            .O(N__13495),
            .I(N__13470));
    InMux I__2404 (
            .O(N__13494),
            .I(N__13465));
    InMux I__2403 (
            .O(N__13491),
            .I(N__13465));
    Span4Mux_s2_v I__2402 (
            .O(N__13488),
            .I(N__13462));
    LocalMux I__2401 (
            .O(N__13483),
            .I(bu_rx_data_3));
    Odrv4 I__2400 (
            .O(N__13478),
            .I(bu_rx_data_3));
    LocalMux I__2399 (
            .O(N__13475),
            .I(bu_rx_data_3));
    Odrv4 I__2398 (
            .O(N__13470),
            .I(bu_rx_data_3));
    LocalMux I__2397 (
            .O(N__13465),
            .I(bu_rx_data_3));
    Odrv4 I__2396 (
            .O(N__13462),
            .I(bu_rx_data_3));
    CEMux I__2395 (
            .O(N__13449),
            .I(N__13422));
    CEMux I__2394 (
            .O(N__13448),
            .I(N__13422));
    CEMux I__2393 (
            .O(N__13447),
            .I(N__13422));
    CEMux I__2392 (
            .O(N__13446),
            .I(N__13422));
    CEMux I__2391 (
            .O(N__13445),
            .I(N__13422));
    CEMux I__2390 (
            .O(N__13444),
            .I(N__13422));
    CEMux I__2389 (
            .O(N__13443),
            .I(N__13422));
    CEMux I__2388 (
            .O(N__13442),
            .I(N__13422));
    CEMux I__2387 (
            .O(N__13441),
            .I(N__13422));
    GlobalMux I__2386 (
            .O(N__13422),
            .I(N__13419));
    gio2CtrlBuf I__2385 (
            .O(N__13419),
            .I(N_76_i_g));
    CascadeMux I__2384 (
            .O(N__13416),
            .I(\buart.Z_rx.bitcountN11_15_i_0_o2_0_cascade_ ));
    InMux I__2383 (
            .O(N__13413),
            .I(N__13408));
    InMux I__2382 (
            .O(N__13412),
            .I(N__13405));
    InMux I__2381 (
            .O(N__13411),
            .I(N__13401));
    LocalMux I__2380 (
            .O(N__13408),
            .I(N__13393));
    LocalMux I__2379 (
            .O(N__13405),
            .I(N__13393));
    InMux I__2378 (
            .O(N__13404),
            .I(N__13390));
    LocalMux I__2377 (
            .O(N__13401),
            .I(N__13387));
    InMux I__2376 (
            .O(N__13400),
            .I(N__13384));
    InMux I__2375 (
            .O(N__13399),
            .I(N__13379));
    InMux I__2374 (
            .O(N__13398),
            .I(N__13379));
    Span4Mux_v I__2373 (
            .O(N__13393),
            .I(N__13376));
    LocalMux I__2372 (
            .O(N__13390),
            .I(N__13373));
    Odrv4 I__2371 (
            .O(N__13387),
            .I(\Lab_UT.scctrl.N_241 ));
    LocalMux I__2370 (
            .O(N__13384),
            .I(\Lab_UT.scctrl.N_241 ));
    LocalMux I__2369 (
            .O(N__13379),
            .I(\Lab_UT.scctrl.N_241 ));
    Odrv4 I__2368 (
            .O(N__13376),
            .I(\Lab_UT.scctrl.N_241 ));
    Odrv4 I__2367 (
            .O(N__13373),
            .I(\Lab_UT.scctrl.N_241 ));
    CascadeMux I__2366 (
            .O(N__13362),
            .I(\Lab_UT.scctrl.g0_70_1_cascade_ ));
    CascadeMux I__2365 (
            .O(N__13359),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0_cascade_ ));
    InMux I__2364 (
            .O(N__13356),
            .I(N__13349));
    InMux I__2363 (
            .O(N__13355),
            .I(N__13349));
    CascadeMux I__2362 (
            .O(N__13354),
            .I(N__13346));
    LocalMux I__2361 (
            .O(N__13349),
            .I(N__13342));
    InMux I__2360 (
            .O(N__13346),
            .I(N__13337));
    InMux I__2359 (
            .O(N__13345),
            .I(N__13337));
    Odrv4 I__2358 (
            .O(N__13342),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0 ));
    LocalMux I__2357 (
            .O(N__13337),
            .I(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0 ));
    InMux I__2356 (
            .O(N__13332),
            .I(N__13329));
    LocalMux I__2355 (
            .O(N__13329),
            .I(buart__rx_shifter_2_fast_6));
    InMux I__2354 (
            .O(N__13326),
            .I(N__13317));
    InMux I__2353 (
            .O(N__13325),
            .I(N__13317));
    InMux I__2352 (
            .O(N__13324),
            .I(N__13317));
    LocalMux I__2351 (
            .O(N__13317),
            .I(\Lab_UT.scctrl.N_444 ));
    CascadeMux I__2350 (
            .O(N__13314),
            .I(N__13310));
    InMux I__2349 (
            .O(N__13313),
            .I(N__13305));
    InMux I__2348 (
            .O(N__13310),
            .I(N__13305));
    LocalMux I__2347 (
            .O(N__13305),
            .I(bu_rx_data_i_2_fast_3));
    InMux I__2346 (
            .O(N__13302),
            .I(N__13299));
    LocalMux I__2345 (
            .O(N__13299),
            .I(N__13296));
    Span4Mux_h I__2344 (
            .O(N__13296),
            .I(N__13293));
    Odrv4 I__2343 (
            .O(N__13293),
            .I(N_243_reti));
    InMux I__2342 (
            .O(N__13290),
            .I(N__13287));
    LocalMux I__2341 (
            .O(N__13287),
            .I(\Lab_UT.scctrl.N_219i ));
    CascadeMux I__2340 (
            .O(N__13284),
            .I(N__13281));
    InMux I__2339 (
            .O(N__13281),
            .I(N__13278));
    LocalMux I__2338 (
            .O(N__13278),
            .I(\Lab_UT.scctrl.N_271_0_0 ));
    CascadeMux I__2337 (
            .O(N__13275),
            .I(\Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_1_cascade_ ));
    InMux I__2336 (
            .O(N__13272),
            .I(N__13269));
    LocalMux I__2335 (
            .O(N__13269),
            .I(\Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0 ));
    CascadeMux I__2334 (
            .O(N__13266),
            .I(\Lab_UT.scctrl.g0_i_o7_1_cascade_ ));
    CascadeMux I__2333 (
            .O(N__13263),
            .I(\Lab_UT.scctrl.N_12_2_cascade_ ));
    InMux I__2332 (
            .O(N__13260),
            .I(N__13255));
    CascadeMux I__2331 (
            .O(N__13259),
            .I(N__13251));
    InMux I__2330 (
            .O(N__13258),
            .I(N__13247));
    LocalMux I__2329 (
            .O(N__13255),
            .I(N__13244));
    InMux I__2328 (
            .O(N__13254),
            .I(N__13241));
    InMux I__2327 (
            .O(N__13251),
            .I(N__13238));
    InMux I__2326 (
            .O(N__13250),
            .I(N__13235));
    LocalMux I__2325 (
            .O(N__13247),
            .I(bu_rx_data_i_2_3_rep1));
    Odrv4 I__2324 (
            .O(N__13244),
            .I(bu_rx_data_i_2_3_rep1));
    LocalMux I__2323 (
            .O(N__13241),
            .I(bu_rx_data_i_2_3_rep1));
    LocalMux I__2322 (
            .O(N__13238),
            .I(bu_rx_data_i_2_3_rep1));
    LocalMux I__2321 (
            .O(N__13235),
            .I(bu_rx_data_i_2_3_rep1));
    CascadeMux I__2320 (
            .O(N__13224),
            .I(N__13220));
    InMux I__2319 (
            .O(N__13223),
            .I(N__13216));
    InMux I__2318 (
            .O(N__13220),
            .I(N__13211));
    InMux I__2317 (
            .O(N__13219),
            .I(N__13211));
    LocalMux I__2316 (
            .O(N__13216),
            .I(N__13208));
    LocalMux I__2315 (
            .O(N__13211),
            .I(N__13205));
    Odrv4 I__2314 (
            .O(N__13208),
            .I(\Lab_UT.scctrl.N_259 ));
    Odrv12 I__2313 (
            .O(N__13205),
            .I(\Lab_UT.scctrl.N_259 ));
    CascadeMux I__2312 (
            .O(N__13200),
            .I(N__13197));
    InMux I__2311 (
            .O(N__13197),
            .I(N__13194));
    LocalMux I__2310 (
            .O(N__13194),
            .I(N__13191));
    Span4Mux_h I__2309 (
            .O(N__13191),
            .I(N__13188));
    Odrv4 I__2308 (
            .O(N__13188),
            .I(\Lab_UT.scctrl.g0_1_i_a8_0_1 ));
    InMux I__2307 (
            .O(N__13185),
            .I(N__13182));
    LocalMux I__2306 (
            .O(N__13182),
            .I(\Lab_UT.scctrl.N_7_0 ));
    InMux I__2305 (
            .O(N__13179),
            .I(N__13176));
    LocalMux I__2304 (
            .O(N__13176),
            .I(\Lab_UT.scctrl.N_10_0 ));
    InMux I__2303 (
            .O(N__13173),
            .I(N__13165));
    InMux I__2302 (
            .O(N__13172),
            .I(N__13165));
    InMux I__2301 (
            .O(N__13171),
            .I(N__13162));
    InMux I__2300 (
            .O(N__13170),
            .I(N__13159));
    LocalMux I__2299 (
            .O(N__13165),
            .I(N__13156));
    LocalMux I__2298 (
            .O(N__13162),
            .I(\Lab_UT.scctrl.N_219 ));
    LocalMux I__2297 (
            .O(N__13159),
            .I(\Lab_UT.scctrl.N_219 ));
    Odrv4 I__2296 (
            .O(N__13156),
            .I(\Lab_UT.scctrl.N_219 ));
    CascadeMux I__2295 (
            .O(N__13149),
            .I(N__13145));
    InMux I__2294 (
            .O(N__13148),
            .I(N__13139));
    InMux I__2293 (
            .O(N__13145),
            .I(N__13139));
    InMux I__2292 (
            .O(N__13144),
            .I(N__13136));
    LocalMux I__2291 (
            .O(N__13139),
            .I(N__13133));
    LocalMux I__2290 (
            .O(N__13136),
            .I(buart__rx_shifter_0_fast_1));
    Odrv4 I__2289 (
            .O(N__13133),
            .I(buart__rx_shifter_0_fast_1));
    InMux I__2288 (
            .O(N__13128),
            .I(N__13125));
    LocalMux I__2287 (
            .O(N__13125),
            .I(\Lab_UT.scctrl.g0_0_i_0 ));
    CascadeMux I__2286 (
            .O(N__13122),
            .I(\Lab_UT.scctrl.g0_0_i_1_cascade_ ));
    CascadeMux I__2285 (
            .O(N__13119),
            .I(\Lab_UT.scctrl.g0_0_i_1_0_cascade_ ));
    InMux I__2284 (
            .O(N__13116),
            .I(N__13113));
    LocalMux I__2283 (
            .O(N__13113),
            .I(\Lab_UT.scctrl.N_5_1 ));
    CascadeMux I__2282 (
            .O(N__13110),
            .I(\Lab_UT.scctrl.g0_2_0_0_a3_1_1_cascade_ ));
    CascadeMux I__2281 (
            .O(N__13107),
            .I(\Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0_cascade_ ));
    InMux I__2280 (
            .O(N__13104),
            .I(N__13101));
    LocalMux I__2279 (
            .O(N__13101),
            .I(\Lab_UT.scctrl.g1_0_5 ));
    CascadeMux I__2278 (
            .O(N__13098),
            .I(\Lab_UT.scctrl.next_state_1_0_2_cascade_ ));
    CascadeMux I__2277 (
            .O(N__13095),
            .I(\Lab_UT.scctrl.N_444_0_cascade_ ));
    InMux I__2276 (
            .O(N__13092),
            .I(N__13089));
    LocalMux I__2275 (
            .O(N__13089),
            .I(\Lab_UT.scctrl.N_319_1_0 ));
    CascadeMux I__2274 (
            .O(N__13086),
            .I(\Lab_UT.scctrl.N_223_1_0_cascade_ ));
    InMux I__2273 (
            .O(N__13083),
            .I(N__13080));
    LocalMux I__2272 (
            .O(N__13080),
            .I(\Lab_UT.scctrl.N_414_1_0 ));
    InMux I__2271 (
            .O(N__13077),
            .I(N__13074));
    LocalMux I__2270 (
            .O(N__13074),
            .I(\Lab_UT.scctrl.N_444_0 ));
    CascadeMux I__2269 (
            .O(N__13071),
            .I(\Lab_UT.scctrl.N_223_1_cascade_ ));
    CascadeMux I__2268 (
            .O(N__13068),
            .I(\Lab_UT.scctrl.N_414_1_cascade_ ));
    InMux I__2267 (
            .O(N__13065),
            .I(N__13062));
    LocalMux I__2266 (
            .O(N__13062),
            .I(N__13058));
    InMux I__2265 (
            .O(N__13061),
            .I(N__13055));
    Odrv4 I__2264 (
            .O(N__13058),
            .I(\Lab_UT.scctrl.g1_0_2_0 ));
    LocalMux I__2263 (
            .O(N__13055),
            .I(\Lab_UT.scctrl.g1_0_2_0 ));
    CascadeMux I__2262 (
            .O(N__13050),
            .I(\Lab_UT.scctrl.next_state_1_2_cascade_ ));
    CascadeMux I__2261 (
            .O(N__13047),
            .I(\Lab_UT.scctrl.N_534_reti_cascade_ ));
    InMux I__2260 (
            .O(N__13044),
            .I(N__13041));
    LocalMux I__2259 (
            .O(N__13041),
            .I(\Lab_UT.scctrl.N_266i ));
    CascadeMux I__2258 (
            .O(N__13038),
            .I(N__13034));
    InMux I__2257 (
            .O(N__13037),
            .I(N__13027));
    InMux I__2256 (
            .O(N__13034),
            .I(N__13024));
    InMux I__2255 (
            .O(N__13033),
            .I(N__13021));
    InMux I__2254 (
            .O(N__13032),
            .I(N__13014));
    InMux I__2253 (
            .O(N__13031),
            .I(N__13011));
    InMux I__2252 (
            .O(N__13030),
            .I(N__13007));
    LocalMux I__2251 (
            .O(N__13027),
            .I(N__13004));
    LocalMux I__2250 (
            .O(N__13024),
            .I(N__13001));
    LocalMux I__2249 (
            .O(N__13021),
            .I(N__12998));
    InMux I__2248 (
            .O(N__13020),
            .I(N__12993));
    InMux I__2247 (
            .O(N__13019),
            .I(N__12993));
    InMux I__2246 (
            .O(N__13018),
            .I(N__12988));
    InMux I__2245 (
            .O(N__13017),
            .I(N__12988));
    LocalMux I__2244 (
            .O(N__13014),
            .I(N__12985));
    LocalMux I__2243 (
            .O(N__13011),
            .I(N__12980));
    InMux I__2242 (
            .O(N__13010),
            .I(N__12977));
    LocalMux I__2241 (
            .O(N__13007),
            .I(N__12971));
    Span12Mux_s7_h I__2240 (
            .O(N__13004),
            .I(N__12968));
    Span4Mux_v I__2239 (
            .O(N__13001),
            .I(N__12957));
    Span4Mux_h I__2238 (
            .O(N__12998),
            .I(N__12957));
    LocalMux I__2237 (
            .O(N__12993),
            .I(N__12957));
    LocalMux I__2236 (
            .O(N__12988),
            .I(N__12957));
    Span4Mux_h I__2235 (
            .O(N__12985),
            .I(N__12957));
    InMux I__2234 (
            .O(N__12984),
            .I(N__12954));
    InMux I__2233 (
            .O(N__12983),
            .I(N__12951));
    Span4Mux_v I__2232 (
            .O(N__12980),
            .I(N__12946));
    LocalMux I__2231 (
            .O(N__12977),
            .I(N__12946));
    InMux I__2230 (
            .O(N__12976),
            .I(N__12939));
    InMux I__2229 (
            .O(N__12975),
            .I(N__12939));
    InMux I__2228 (
            .O(N__12974),
            .I(N__12939));
    Odrv4 I__2227 (
            .O(N__12971),
            .I(bu_rx_data_2));
    Odrv12 I__2226 (
            .O(N__12968),
            .I(bu_rx_data_2));
    Odrv4 I__2225 (
            .O(N__12957),
            .I(bu_rx_data_2));
    LocalMux I__2224 (
            .O(N__12954),
            .I(bu_rx_data_2));
    LocalMux I__2223 (
            .O(N__12951),
            .I(bu_rx_data_2));
    Odrv4 I__2222 (
            .O(N__12946),
            .I(bu_rx_data_2));
    LocalMux I__2221 (
            .O(N__12939),
            .I(bu_rx_data_2));
    CascadeMux I__2220 (
            .O(N__12924),
            .I(N__12921));
    InMux I__2219 (
            .O(N__12921),
            .I(N__12918));
    LocalMux I__2218 (
            .O(N__12918),
            .I(N__12915));
    Span4Mux_v I__2217 (
            .O(N__12915),
            .I(N__12911));
    InMux I__2216 (
            .O(N__12914),
            .I(N__12908));
    Odrv4 I__2215 (
            .O(N__12911),
            .I(\Lab_UT.N_540 ));
    LocalMux I__2214 (
            .O(N__12908),
            .I(\Lab_UT.N_540 ));
    InMux I__2213 (
            .O(N__12903),
            .I(N__12900));
    LocalMux I__2212 (
            .O(N__12900),
            .I(\Lab_UT.scctrl.N_399_0 ));
    InMux I__2211 (
            .O(N__12897),
            .I(N__12894));
    LocalMux I__2210 (
            .O(N__12894),
            .I(\Lab_UT.scctrl.sccEldByte_i_a2_0Z0Z_1 ));
    InMux I__2209 (
            .O(N__12891),
            .I(N__12888));
    LocalMux I__2208 (
            .O(N__12888),
            .I(\Lab_UT.scctrl.g2 ));
    InMux I__2207 (
            .O(N__12885),
            .I(N__12882));
    LocalMux I__2206 (
            .O(N__12882),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18 ));
    InMux I__2205 (
            .O(N__12879),
            .I(N__12875));
    CascadeMux I__2204 (
            .O(N__12878),
            .I(N__12872));
    LocalMux I__2203 (
            .O(N__12875),
            .I(N__12869));
    InMux I__2202 (
            .O(N__12872),
            .I(N__12866));
    Odrv4 I__2201 (
            .O(N__12869),
            .I(\Lab_UT.scdp.key0_4 ));
    LocalMux I__2200 (
            .O(N__12866),
            .I(\Lab_UT.scdp.key0_4 ));
    InMux I__2199 (
            .O(N__12861),
            .I(N__12855));
    InMux I__2198 (
            .O(N__12860),
            .I(N__12855));
    LocalMux I__2197 (
            .O(N__12855),
            .I(\Lab_UT.scdp.prng_lfsr_4 ));
    InMux I__2196 (
            .O(N__12852),
            .I(N__12849));
    LocalMux I__2195 (
            .O(N__12849),
            .I(N__12845));
    InMux I__2194 (
            .O(N__12848),
            .I(N__12842));
    Odrv4 I__2193 (
            .O(N__12845),
            .I(\Lab_UT.scdp.key3_4 ));
    LocalMux I__2192 (
            .O(N__12842),
            .I(\Lab_UT.scdp.key3_4 ));
    InMux I__2191 (
            .O(N__12837),
            .I(N__12834));
    LocalMux I__2190 (
            .O(N__12834),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28 ));
    InMux I__2189 (
            .O(N__12831),
            .I(N__12825));
    InMux I__2188 (
            .O(N__12830),
            .I(N__12825));
    LocalMux I__2187 (
            .O(N__12825),
            .I(N__12822));
    Span4Mux_h I__2186 (
            .O(N__12822),
            .I(N__12819));
    Odrv4 I__2185 (
            .O(N__12819),
            .I(\Lab_UT.scdp.prng_lfsr_11 ));
    CascadeMux I__2184 (
            .O(N__12816),
            .I(N__12813));
    InMux I__2183 (
            .O(N__12813),
            .I(N__12810));
    LocalMux I__2182 (
            .O(N__12810),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26 ));
    InMux I__2181 (
            .O(N__12807),
            .I(N__12801));
    InMux I__2180 (
            .O(N__12806),
            .I(N__12801));
    LocalMux I__2179 (
            .O(N__12801),
            .I(\Lab_UT.scdp.prng_lfsr_12 ));
    InMux I__2178 (
            .O(N__12798),
            .I(N__12795));
    LocalMux I__2177 (
            .O(N__12795),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9 ));
    CEMux I__2176 (
            .O(N__12792),
            .I(N__12765));
    CEMux I__2175 (
            .O(N__12791),
            .I(N__12765));
    CEMux I__2174 (
            .O(N__12790),
            .I(N__12765));
    CEMux I__2173 (
            .O(N__12789),
            .I(N__12765));
    CEMux I__2172 (
            .O(N__12788),
            .I(N__12765));
    CEMux I__2171 (
            .O(N__12787),
            .I(N__12765));
    CEMux I__2170 (
            .O(N__12786),
            .I(N__12765));
    CEMux I__2169 (
            .O(N__12785),
            .I(N__12765));
    CEMux I__2168 (
            .O(N__12784),
            .I(N__12765));
    GlobalMux I__2167 (
            .O(N__12765),
            .I(N__12762));
    gio2CtrlBuf I__2166 (
            .O(N__12762),
            .I(\Lab_UT.sccLdLFSR_g ));
    InMux I__2165 (
            .O(N__12759),
            .I(N__12756));
    LocalMux I__2164 (
            .O(N__12756),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16 ));
    CascadeMux I__2163 (
            .O(N__12753),
            .I(N__12750));
    InMux I__2162 (
            .O(N__12750),
            .I(N__12747));
    LocalMux I__2161 (
            .O(N__12747),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24 ));
    InMux I__2160 (
            .O(N__12744),
            .I(N__12741));
    LocalMux I__2159 (
            .O(N__12741),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0 ));
    CascadeMux I__2158 (
            .O(N__12738),
            .I(\Lab_UT.scdp.d2eData_3_0_cascade_ ));
    InMux I__2157 (
            .O(N__12735),
            .I(N__12732));
    LocalMux I__2156 (
            .O(N__12732),
            .I(N__12729));
    Span4Mux_h I__2155 (
            .O(N__12729),
            .I(N__12725));
    InMux I__2154 (
            .O(N__12728),
            .I(N__12722));
    Odrv4 I__2153 (
            .O(N__12725),
            .I(\Lab_UT.scdp.N_262_i ));
    LocalMux I__2152 (
            .O(N__12722),
            .I(\Lab_UT.scdp.N_262_i ));
    InMux I__2151 (
            .O(N__12717),
            .I(N__12714));
    LocalMux I__2150 (
            .O(N__12714),
            .I(N__12711));
    Odrv12 I__2149 (
            .O(N__12711),
            .I(\Lab_UT.scdp.u1.g0_0_i_a5_0_0 ));
    InMux I__2148 (
            .O(N__12708),
            .I(N__12702));
    InMux I__2147 (
            .O(N__12707),
            .I(N__12702));
    LocalMux I__2146 (
            .O(N__12702),
            .I(N__12699));
    Span4Mux_h I__2145 (
            .O(N__12699),
            .I(N__12695));
    InMux I__2144 (
            .O(N__12698),
            .I(N__12692));
    Span4Mux_v I__2143 (
            .O(N__12695),
            .I(N__12687));
    LocalMux I__2142 (
            .O(N__12692),
            .I(N__12684));
    InMux I__2141 (
            .O(N__12691),
            .I(N__12679));
    InMux I__2140 (
            .O(N__12690),
            .I(N__12679));
    Odrv4 I__2139 (
            .O(N__12687),
            .I(\Lab_UT.scdp.d2eData_3_0 ));
    Odrv4 I__2138 (
            .O(N__12684),
            .I(\Lab_UT.scdp.d2eData_3_0 ));
    LocalMux I__2137 (
            .O(N__12679),
            .I(\Lab_UT.scdp.d2eData_3_0 ));
    CascadeMux I__2136 (
            .O(N__12672),
            .I(N__12668));
    InMux I__2135 (
            .O(N__12671),
            .I(N__12660));
    InMux I__2134 (
            .O(N__12668),
            .I(N__12660));
    InMux I__2133 (
            .O(N__12667),
            .I(N__12655));
    InMux I__2132 (
            .O(N__12666),
            .I(N__12655));
    InMux I__2131 (
            .O(N__12665),
            .I(N__12652));
    LocalMux I__2130 (
            .O(N__12660),
            .I(N__12649));
    LocalMux I__2129 (
            .O(N__12655),
            .I(N__12646));
    LocalMux I__2128 (
            .O(N__12652),
            .I(\Lab_UT.scdp.u1.byteToDecryptZ0Z_2 ));
    Odrv4 I__2127 (
            .O(N__12649),
            .I(\Lab_UT.scdp.u1.byteToDecryptZ0Z_2 ));
    Odrv12 I__2126 (
            .O(N__12646),
            .I(\Lab_UT.scdp.u1.byteToDecryptZ0Z_2 ));
    InMux I__2125 (
            .O(N__12639),
            .I(N__12627));
    InMux I__2124 (
            .O(N__12638),
            .I(N__12627));
    InMux I__2123 (
            .O(N__12637),
            .I(N__12627));
    InMux I__2122 (
            .O(N__12636),
            .I(N__12627));
    LocalMux I__2121 (
            .O(N__12627),
            .I(N__12622));
    InMux I__2120 (
            .O(N__12626),
            .I(N__12617));
    InMux I__2119 (
            .O(N__12625),
            .I(N__12617));
    Span12Mux_s4_h I__2118 (
            .O(N__12622),
            .I(N__12613));
    LocalMux I__2117 (
            .O(N__12617),
            .I(N__12610));
    InMux I__2116 (
            .O(N__12616),
            .I(N__12607));
    Odrv12 I__2115 (
            .O(N__12613),
            .I(\Lab_UT.scdp.d2eData_3_2 ));
    Odrv4 I__2114 (
            .O(N__12610),
            .I(\Lab_UT.scdp.d2eData_3_2 ));
    LocalMux I__2113 (
            .O(N__12607),
            .I(\Lab_UT.scdp.d2eData_3_2 ));
    InMux I__2112 (
            .O(N__12600),
            .I(N__12597));
    LocalMux I__2111 (
            .O(N__12597),
            .I(N__12594));
    Odrv4 I__2110 (
            .O(N__12594),
            .I(\Lab_UT.scdp.u1.g0_0_i_a5_0_0_0 ));
    InMux I__2109 (
            .O(N__12591),
            .I(N__12588));
    LocalMux I__2108 (
            .O(N__12588),
            .I(N__12584));
    CascadeMux I__2107 (
            .O(N__12587),
            .I(N__12581));
    Span4Mux_v I__2106 (
            .O(N__12584),
            .I(N__12578));
    InMux I__2105 (
            .O(N__12581),
            .I(N__12575));
    Odrv4 I__2104 (
            .O(N__12578),
            .I(\Lab_UT.scdp.key0_6 ));
    LocalMux I__2103 (
            .O(N__12575),
            .I(\Lab_UT.scdp.key0_6 ));
    InMux I__2102 (
            .O(N__12570),
            .I(N__12565));
    InMux I__2101 (
            .O(N__12569),
            .I(N__12560));
    InMux I__2100 (
            .O(N__12568),
            .I(N__12560));
    LocalMux I__2099 (
            .O(N__12565),
            .I(N__12557));
    LocalMux I__2098 (
            .O(N__12560),
            .I(N__12554));
    Span4Mux_h I__2097 (
            .O(N__12557),
            .I(N__12551));
    Span4Mux_h I__2096 (
            .O(N__12554),
            .I(N__12548));
    Odrv4 I__2095 (
            .O(N__12551),
            .I(\Lab_UT.scdp.prng_lfsr_6 ));
    Odrv4 I__2094 (
            .O(N__12548),
            .I(\Lab_UT.scdp.prng_lfsr_6 ));
    InMux I__2093 (
            .O(N__12543),
            .I(N__12540));
    LocalMux I__2092 (
            .O(N__12540),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20 ));
    InMux I__2091 (
            .O(N__12537),
            .I(N__12534));
    LocalMux I__2090 (
            .O(N__12534),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8 ));
    CascadeMux I__2089 (
            .O(N__12531),
            .I(\Lab_UT.scctrl.N_22_i_cascade_ ));
    CascadeMux I__2088 (
            .O(N__12528),
            .I(\Lab_UT.state_1_ret_0_RNI9C1NH_0_cascade_ ));
    InMux I__2087 (
            .O(N__12525),
            .I(N__12521));
    InMux I__2086 (
            .O(N__12524),
            .I(N__12518));
    LocalMux I__2085 (
            .O(N__12521),
            .I(\Lab_UT.scdp.key3_5 ));
    LocalMux I__2084 (
            .O(N__12518),
            .I(\Lab_UT.scdp.key3_5 ));
    InMux I__2083 (
            .O(N__12513),
            .I(N__12504));
    InMux I__2082 (
            .O(N__12512),
            .I(N__12504));
    InMux I__2081 (
            .O(N__12511),
            .I(N__12504));
    LocalMux I__2080 (
            .O(N__12504),
            .I(\Lab_UT.state_1_ret_0_RNI9C1NH_0 ));
    InMux I__2079 (
            .O(N__12501),
            .I(N__12498));
    LocalMux I__2078 (
            .O(N__12498),
            .I(N__12494));
    CascadeMux I__2077 (
            .O(N__12497),
            .I(N__12491));
    Span4Mux_v I__2076 (
            .O(N__12494),
            .I(N__12488));
    InMux I__2075 (
            .O(N__12491),
            .I(N__12485));
    Odrv4 I__2074 (
            .O(N__12488),
            .I(\Lab_UT.scdp.key3_6 ));
    LocalMux I__2073 (
            .O(N__12485),
            .I(\Lab_UT.scdp.key3_6 ));
    InMux I__2072 (
            .O(N__12480),
            .I(N__12473));
    InMux I__2071 (
            .O(N__12479),
            .I(N__12468));
    InMux I__2070 (
            .O(N__12478),
            .I(N__12468));
    InMux I__2069 (
            .O(N__12477),
            .I(N__12463));
    InMux I__2068 (
            .O(N__12476),
            .I(N__12463));
    LocalMux I__2067 (
            .O(N__12473),
            .I(\Lab_UT.state_1_RNI6EDGH_0_2 ));
    LocalMux I__2066 (
            .O(N__12468),
            .I(\Lab_UT.state_1_RNI6EDGH_0_2 ));
    LocalMux I__2065 (
            .O(N__12463),
            .I(\Lab_UT.state_1_RNI6EDGH_0_2 ));
    CascadeMux I__2064 (
            .O(N__12456),
            .I(N__12452));
    InMux I__2063 (
            .O(N__12455),
            .I(N__12449));
    InMux I__2062 (
            .O(N__12452),
            .I(N__12446));
    LocalMux I__2061 (
            .O(N__12449),
            .I(\Lab_UT.scdp.key0_5 ));
    LocalMux I__2060 (
            .O(N__12446),
            .I(\Lab_UT.scdp.key0_5 ));
    InMux I__2059 (
            .O(N__12441),
            .I(N__12438));
    LocalMux I__2058 (
            .O(N__12438),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    InMux I__2057 (
            .O(N__12435),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__2056 (
            .O(N__12432),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    CEMux I__2055 (
            .O(N__12429),
            .I(N__12426));
    LocalMux I__2054 (
            .O(N__12426),
            .I(N__12422));
    CEMux I__2053 (
            .O(N__12425),
            .I(N__12419));
    Span4Mux_v I__2052 (
            .O(N__12422),
            .I(N__12416));
    LocalMux I__2051 (
            .O(N__12419),
            .I(N__12413));
    Span4Mux_h I__2050 (
            .O(N__12416),
            .I(N__12410));
    Sp12to4 I__2049 (
            .O(N__12413),
            .I(N__12407));
    Odrv4 I__2048 (
            .O(N__12410),
            .I(\buart.Z_rx.N_78 ));
    Odrv12 I__2047 (
            .O(N__12407),
            .I(\buart.Z_rx.N_78 ));
    CascadeMux I__2046 (
            .O(N__12402),
            .I(\Lab_UT.scctrl.N_418_0_cascade_ ));
    InMux I__2045 (
            .O(N__12399),
            .I(N__12396));
    LocalMux I__2044 (
            .O(N__12396),
            .I(\Lab_UT.scctrl.g0_2 ));
    CascadeMux I__2043 (
            .O(N__12393),
            .I(\Lab_UT.scctrl.g0_2_cascade_ ));
    InMux I__2042 (
            .O(N__12390),
            .I(N__12384));
    InMux I__2041 (
            .O(N__12389),
            .I(N__12384));
    LocalMux I__2040 (
            .O(N__12384),
            .I(N__12381));
    Odrv4 I__2039 (
            .O(N__12381),
            .I(\Lab_UT.scctrl.g1_1 ));
    CascadeMux I__2038 (
            .O(N__12378),
            .I(\Lab_UT.scctrl.N_418_2_0_cascade_ ));
    InMux I__2037 (
            .O(N__12375),
            .I(N__12372));
    LocalMux I__2036 (
            .O(N__12372),
            .I(N__12369));
    Span12Mux_s3_v I__2035 (
            .O(N__12369),
            .I(N__12366));
    Odrv12 I__2034 (
            .O(N__12366),
            .I(\Lab_UT.scctrl.g1_1_2 ));
    CascadeMux I__2033 (
            .O(N__12363),
            .I(\Lab_UT.scctrl.N_39_i_cascade_ ));
    CascadeMux I__2032 (
            .O(N__12360),
            .I(CONSTANT_ONE_NET_cascade_));
    InMux I__2031 (
            .O(N__12357),
            .I(N__12354));
    LocalMux I__2030 (
            .O(N__12354),
            .I(N__12351));
    Span4Mux_v I__2029 (
            .O(N__12351),
            .I(N__12348));
    Odrv4 I__2028 (
            .O(N__12348),
            .I(\ufifo.sb_ram512x8_inst_RNIKTQ21 ));
    InMux I__2027 (
            .O(N__12345),
            .I(N__12342));
    LocalMux I__2026 (
            .O(N__12342),
            .I(N__12339));
    Span4Mux_v I__2025 (
            .O(N__12339),
            .I(N__12336));
    Span4Mux_h I__2024 (
            .O(N__12336),
            .I(N__12333));
    Odrv4 I__2023 (
            .O(N__12333),
            .I(\ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1Z0Z_0 ));
    InMux I__2022 (
            .O(N__12330),
            .I(N__12327));
    LocalMux I__2021 (
            .O(N__12327),
            .I(N__12317));
    InMux I__2020 (
            .O(N__12326),
            .I(N__12299));
    InMux I__2019 (
            .O(N__12325),
            .I(N__12299));
    InMux I__2018 (
            .O(N__12324),
            .I(N__12299));
    InMux I__2017 (
            .O(N__12323),
            .I(N__12299));
    InMux I__2016 (
            .O(N__12322),
            .I(N__12299));
    InMux I__2015 (
            .O(N__12321),
            .I(N__12294));
    InMux I__2014 (
            .O(N__12320),
            .I(N__12294));
    Span4Mux_v I__2013 (
            .O(N__12317),
            .I(N__12291));
    InMux I__2012 (
            .O(N__12316),
            .I(N__12288));
    InMux I__2011 (
            .O(N__12315),
            .I(N__12281));
    InMux I__2010 (
            .O(N__12314),
            .I(N__12281));
    InMux I__2009 (
            .O(N__12313),
            .I(N__12281));
    InMux I__2008 (
            .O(N__12312),
            .I(N__12274));
    InMux I__2007 (
            .O(N__12311),
            .I(N__12274));
    InMux I__2006 (
            .O(N__12310),
            .I(N__12274));
    LocalMux I__2005 (
            .O(N__12299),
            .I(N__12269));
    LocalMux I__2004 (
            .O(N__12294),
            .I(N__12269));
    Span4Mux_h I__2003 (
            .O(N__12291),
            .I(N__12264));
    LocalMux I__2002 (
            .O(N__12288),
            .I(N__12264));
    LocalMux I__2001 (
            .O(N__12281),
            .I(N_368));
    LocalMux I__2000 (
            .O(N__12274),
            .I(N_368));
    Odrv4 I__1999 (
            .O(N__12269),
            .I(N_368));
    Odrv4 I__1998 (
            .O(N__12264),
            .I(N_368));
    InMux I__1997 (
            .O(N__12255),
            .I(N__12252));
    LocalMux I__1996 (
            .O(N__12252),
            .I(N__12249));
    Span4Mux_h I__1995 (
            .O(N__12249),
            .I(N__12246));
    Span4Mux_v I__1994 (
            .O(N__12246),
            .I(N__12243));
    Odrv4 I__1993 (
            .O(N__12243),
            .I(utb_txdata_0));
    CascadeMux I__1992 (
            .O(N__12240),
            .I(N__12237));
    InMux I__1991 (
            .O(N__12237),
            .I(N__12234));
    LocalMux I__1990 (
            .O(N__12234),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    InMux I__1989 (
            .O(N__12231),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    CascadeMux I__1988 (
            .O(N__12228),
            .I(N__12225));
    InMux I__1987 (
            .O(N__12225),
            .I(N__12222));
    LocalMux I__1986 (
            .O(N__12222),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__1985 (
            .O(N__12219),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    InMux I__1984 (
            .O(N__12216),
            .I(N__12213));
    LocalMux I__1983 (
            .O(N__12213),
            .I(N__12210));
    Odrv4 I__1982 (
            .O(N__12210),
            .I(\Lab_UT.scctrl.N_263_0 ));
    InMux I__1981 (
            .O(N__12207),
            .I(N__12204));
    LocalMux I__1980 (
            .O(N__12204),
            .I(\Lab_UT.scctrl.N_233_0 ));
    InMux I__1979 (
            .O(N__12201),
            .I(N__12198));
    LocalMux I__1978 (
            .O(N__12198),
            .I(\Lab_UT.scctrl.N_351_1_0 ));
    CascadeMux I__1977 (
            .O(N__12195),
            .I(\Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_5_1_cascade_ ));
    CascadeMux I__1976 (
            .O(N__12192),
            .I(N__12189));
    InMux I__1975 (
            .O(N__12189),
            .I(N__12185));
    CascadeMux I__1974 (
            .O(N__12188),
            .I(N__12182));
    LocalMux I__1973 (
            .O(N__12185),
            .I(N__12179));
    InMux I__1972 (
            .O(N__12182),
            .I(N__12176));
    Odrv4 I__1971 (
            .O(N__12179),
            .I(\Lab_UT.N_540i ));
    LocalMux I__1970 (
            .O(N__12176),
            .I(\Lab_UT.N_540i ));
    InMux I__1969 (
            .O(N__12171),
            .I(N__12168));
    LocalMux I__1968 (
            .O(N__12168),
            .I(\Lab_UT.scctrl.N_266 ));
    InMux I__1967 (
            .O(N__12165),
            .I(N__12161));
    InMux I__1966 (
            .O(N__12164),
            .I(N__12158));
    LocalMux I__1965 (
            .O(N__12161),
            .I(N__12155));
    LocalMux I__1964 (
            .O(N__12158),
            .I(\Lab_UT.scctrl.N_472_0 ));
    Odrv12 I__1963 (
            .O(N__12155),
            .I(\Lab_UT.scctrl.N_472_0 ));
    InMux I__1962 (
            .O(N__12150),
            .I(N__12147));
    LocalMux I__1961 (
            .O(N__12147),
            .I(\Lab_UT.scctrl.N_241_reti ));
    CascadeMux I__1960 (
            .O(N__12144),
            .I(\Lab_UT.scctrl.N_241_reti_cascade_ ));
    CascadeMux I__1959 (
            .O(N__12141),
            .I(N__12138));
    InMux I__1958 (
            .O(N__12138),
            .I(N__12135));
    LocalMux I__1957 (
            .O(N__12135),
            .I(N__12132));
    Odrv4 I__1956 (
            .O(N__12132),
            .I(\Lab_UT.scctrl.N_319_0 ));
    InMux I__1955 (
            .O(N__12129),
            .I(N__12126));
    LocalMux I__1954 (
            .O(N__12126),
            .I(N__12123));
    Odrv4 I__1953 (
            .O(N__12123),
            .I(\Lab_UT.scctrl.N_414_0 ));
    CascadeMux I__1952 (
            .O(N__12120),
            .I(\Lab_UT.scctrl.N_415_1_cascade_ ));
    InMux I__1951 (
            .O(N__12117),
            .I(N__12114));
    LocalMux I__1950 (
            .O(N__12114),
            .I(\Lab_UT.scctrl.g1_0_0_0 ));
    InMux I__1949 (
            .O(N__12111),
            .I(N__12108));
    LocalMux I__1948 (
            .O(N__12108),
            .I(\Lab_UT.scctrl.N_259i ));
    InMux I__1947 (
            .O(N__12105),
            .I(N__12102));
    LocalMux I__1946 (
            .O(N__12102),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10 ));
    InMux I__1945 (
            .O(N__12099),
            .I(N__12096));
    LocalMux I__1944 (
            .O(N__12096),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2 ));
    CascadeMux I__1943 (
            .O(N__12093),
            .I(\Lab_UT.scdp.d2eData_3_2_cascade_ ));
    InMux I__1942 (
            .O(N__12090),
            .I(N__12085));
    InMux I__1941 (
            .O(N__12089),
            .I(N__12082));
    InMux I__1940 (
            .O(N__12088),
            .I(N__12078));
    LocalMux I__1939 (
            .O(N__12085),
            .I(N__12073));
    LocalMux I__1938 (
            .O(N__12082),
            .I(N__12073));
    InMux I__1937 (
            .O(N__12081),
            .I(N__12070));
    LocalMux I__1936 (
            .O(N__12078),
            .I(N__12067));
    Span4Mux_v I__1935 (
            .O(N__12073),
            .I(N__12064));
    LocalMux I__1934 (
            .O(N__12070),
            .I(N__12061));
    Span4Mux_v I__1933 (
            .O(N__12067),
            .I(N__12056));
    Span4Mux_h I__1932 (
            .O(N__12064),
            .I(N__12056));
    Span4Mux_h I__1931 (
            .O(N__12061),
            .I(N__12053));
    Odrv4 I__1930 (
            .O(N__12056),
            .I(\Lab_UT.scdp.N_234_i ));
    Odrv4 I__1929 (
            .O(N__12053),
            .I(\Lab_UT.scdp.N_234_i ));
    CascadeMux I__1928 (
            .O(N__12048),
            .I(N__12044));
    InMux I__1927 (
            .O(N__12047),
            .I(N__12040));
    InMux I__1926 (
            .O(N__12044),
            .I(N__12037));
    CascadeMux I__1925 (
            .O(N__12043),
            .I(N__12031));
    LocalMux I__1924 (
            .O(N__12040),
            .I(N__12026));
    LocalMux I__1923 (
            .O(N__12037),
            .I(N__12026));
    InMux I__1922 (
            .O(N__12036),
            .I(N__12023));
    InMux I__1921 (
            .O(N__12035),
            .I(N__12018));
    InMux I__1920 (
            .O(N__12034),
            .I(N__12015));
    InMux I__1919 (
            .O(N__12031),
            .I(N__12012));
    Sp12to4 I__1918 (
            .O(N__12026),
            .I(N__12007));
    LocalMux I__1917 (
            .O(N__12023),
            .I(N__12007));
    InMux I__1916 (
            .O(N__12022),
            .I(N__12004));
    InMux I__1915 (
            .O(N__12021),
            .I(N__12001));
    LocalMux I__1914 (
            .O(N__12018),
            .I(\Lab_UT.scdp.byteToDecrypt_5 ));
    LocalMux I__1913 (
            .O(N__12015),
            .I(\Lab_UT.scdp.byteToDecrypt_5 ));
    LocalMux I__1912 (
            .O(N__12012),
            .I(\Lab_UT.scdp.byteToDecrypt_5 ));
    Odrv12 I__1911 (
            .O(N__12007),
            .I(\Lab_UT.scdp.byteToDecrypt_5 ));
    LocalMux I__1910 (
            .O(N__12004),
            .I(\Lab_UT.scdp.byteToDecrypt_5 ));
    LocalMux I__1909 (
            .O(N__12001),
            .I(\Lab_UT.scdp.byteToDecrypt_5 ));
    InMux I__1908 (
            .O(N__11988),
            .I(N__11985));
    LocalMux I__1907 (
            .O(N__11985),
            .I(N__11982));
    Odrv4 I__1906 (
            .O(N__11982),
            .I(\Lab_UT.scdp.N_228_i_0 ));
    CascadeMux I__1905 (
            .O(N__11979),
            .I(\Lab_UT.scdp.g0_0_i_0_cascade_ ));
    InMux I__1904 (
            .O(N__11976),
            .I(N__11964));
    InMux I__1903 (
            .O(N__11975),
            .I(N__11964));
    InMux I__1902 (
            .O(N__11974),
            .I(N__11964));
    InMux I__1901 (
            .O(N__11973),
            .I(N__11959));
    InMux I__1900 (
            .O(N__11972),
            .I(N__11956));
    InMux I__1899 (
            .O(N__11971),
            .I(N__11952));
    LocalMux I__1898 (
            .O(N__11964),
            .I(N__11949));
    InMux I__1897 (
            .O(N__11963),
            .I(N__11946));
    InMux I__1896 (
            .O(N__11962),
            .I(N__11943));
    LocalMux I__1895 (
            .O(N__11959),
            .I(N__11938));
    LocalMux I__1894 (
            .O(N__11956),
            .I(N__11938));
    InMux I__1893 (
            .O(N__11955),
            .I(N__11935));
    LocalMux I__1892 (
            .O(N__11952),
            .I(\Lab_UT.scdp.d2eData_3_5 ));
    Odrv4 I__1891 (
            .O(N__11949),
            .I(\Lab_UT.scdp.d2eData_3_5 ));
    LocalMux I__1890 (
            .O(N__11946),
            .I(\Lab_UT.scdp.d2eData_3_5 ));
    LocalMux I__1889 (
            .O(N__11943),
            .I(\Lab_UT.scdp.d2eData_3_5 ));
    Odrv4 I__1888 (
            .O(N__11938),
            .I(\Lab_UT.scdp.d2eData_3_5 ));
    LocalMux I__1887 (
            .O(N__11935),
            .I(\Lab_UT.scdp.d2eData_3_5 ));
    InMux I__1886 (
            .O(N__11922),
            .I(N__11919));
    LocalMux I__1885 (
            .O(N__11919),
            .I(N__11916));
    Span4Mux_h I__1884 (
            .O(N__11916),
            .I(N__11913));
    Odrv4 I__1883 (
            .O(N__11913),
            .I(\Lab_UT.scdp.g0_0_i_1_1 ));
    CascadeMux I__1882 (
            .O(N__11910),
            .I(\Lab_UT.scctrl.g1_1_1_1_cascade_ ));
    InMux I__1881 (
            .O(N__11907),
            .I(N__11904));
    LocalMux I__1880 (
            .O(N__11904),
            .I(\Lab_UT.scctrl.g2_0 ));
    CascadeMux I__1879 (
            .O(N__11901),
            .I(N__11898));
    InMux I__1878 (
            .O(N__11898),
            .I(N__11895));
    LocalMux I__1877 (
            .O(N__11895),
            .I(\Lab_UT.scctrl.g1_3 ));
    InMux I__1876 (
            .O(N__11892),
            .I(N__11889));
    LocalMux I__1875 (
            .O(N__11889),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27 ));
    CascadeMux I__1874 (
            .O(N__11886),
            .I(N__11883));
    InMux I__1873 (
            .O(N__11883),
            .I(N__11880));
    LocalMux I__1872 (
            .O(N__11880),
            .I(N__11877));
    Span4Mux_h I__1871 (
            .O(N__11877),
            .I(N__11874));
    Odrv4 I__1870 (
            .O(N__11874),
            .I(\Lab_UT.scdp.byteToEncrypt_4 ));
    InMux I__1869 (
            .O(N__11871),
            .I(N__11862));
    InMux I__1868 (
            .O(N__11870),
            .I(N__11862));
    InMux I__1867 (
            .O(N__11869),
            .I(N__11862));
    LocalMux I__1866 (
            .O(N__11862),
            .I(N__11859));
    Span4Mux_h I__1865 (
            .O(N__11859),
            .I(N__11856));
    Odrv4 I__1864 (
            .O(N__11856),
            .I(\Lab_UT.scdp.b2a0.N_258_i ));
    InMux I__1863 (
            .O(N__11853),
            .I(N__11850));
    LocalMux I__1862 (
            .O(N__11850),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1 ));
    InMux I__1861 (
            .O(N__11847),
            .I(N__11842));
    InMux I__1860 (
            .O(N__11846),
            .I(N__11837));
    InMux I__1859 (
            .O(N__11845),
            .I(N__11834));
    LocalMux I__1858 (
            .O(N__11842),
            .I(N__11831));
    InMux I__1857 (
            .O(N__11841),
            .I(N__11827));
    InMux I__1856 (
            .O(N__11840),
            .I(N__11824));
    LocalMux I__1855 (
            .O(N__11837),
            .I(N__11817));
    LocalMux I__1854 (
            .O(N__11834),
            .I(N__11817));
    Span4Mux_v I__1853 (
            .O(N__11831),
            .I(N__11817));
    InMux I__1852 (
            .O(N__11830),
            .I(N__11814));
    LocalMux I__1851 (
            .O(N__11827),
            .I(\Lab_UT.scdp.d2eData_3_1_1 ));
    LocalMux I__1850 (
            .O(N__11824),
            .I(\Lab_UT.scdp.d2eData_3_1_1 ));
    Odrv4 I__1849 (
            .O(N__11817),
            .I(\Lab_UT.scdp.d2eData_3_1_1 ));
    LocalMux I__1848 (
            .O(N__11814),
            .I(\Lab_UT.scdp.d2eData_3_1_1 ));
    InMux I__1847 (
            .O(N__11805),
            .I(N__11802));
    LocalMux I__1846 (
            .O(N__11802),
            .I(\Lab_UT.scdp.d2eData_3_0_a2_0_4 ));
    CascadeMux I__1845 (
            .O(N__11799),
            .I(\Lab_UT.scdp.d2eData_3_0_a2_0_4_cascade_ ));
    InMux I__1844 (
            .O(N__11796),
            .I(N__11793));
    LocalMux I__1843 (
            .O(N__11793),
            .I(N__11788));
    InMux I__1842 (
            .O(N__11792),
            .I(N__11783));
    InMux I__1841 (
            .O(N__11791),
            .I(N__11783));
    Odrv4 I__1840 (
            .O(N__11788),
            .I(\Lab_UT.scdp.N_246_i ));
    LocalMux I__1839 (
            .O(N__11783),
            .I(\Lab_UT.scdp.N_246_i ));
    CascadeMux I__1838 (
            .O(N__11778),
            .I(\Lab_UT.scdp.N_246_i_cascade_ ));
    InMux I__1837 (
            .O(N__11775),
            .I(N__11772));
    LocalMux I__1836 (
            .O(N__11772),
            .I(\Lab_UT.scdp.u0.L4_tx_data_0_a2_1_6 ));
    InMux I__1835 (
            .O(N__11769),
            .I(N__11766));
    LocalMux I__1834 (
            .O(N__11766),
            .I(\Lab_UT.scdp.N_256_i ));
    InMux I__1833 (
            .O(N__11763),
            .I(N__11759));
    CascadeMux I__1832 (
            .O(N__11762),
            .I(N__11756));
    LocalMux I__1831 (
            .O(N__11759),
            .I(N__11753));
    InMux I__1830 (
            .O(N__11756),
            .I(N__11750));
    Odrv12 I__1829 (
            .O(N__11753),
            .I(\Lab_UT.scdp.key0_2 ));
    LocalMux I__1828 (
            .O(N__11750),
            .I(\Lab_UT.scdp.key0_2 ));
    CascadeMux I__1827 (
            .O(N__11745),
            .I(\Lab_UT.scdp.u1.g0_0_i_a5_0_0_1_cascade_ ));
    InMux I__1826 (
            .O(N__11742),
            .I(N__11739));
    LocalMux I__1825 (
            .O(N__11739),
            .I(\Lab_UT.scdp.u1.g0_0_i_a5_0_2_1 ));
    InMux I__1824 (
            .O(N__11736),
            .I(N__11733));
    LocalMux I__1823 (
            .O(N__11733),
            .I(\Lab_UT.scdp.N_6_1 ));
    CascadeMux I__1822 (
            .O(N__11730),
            .I(\Lab_UT.scdp.d2eData_3_0_3_cascade_ ));
    InMux I__1821 (
            .O(N__11727),
            .I(N__11721));
    InMux I__1820 (
            .O(N__11726),
            .I(N__11721));
    LocalMux I__1819 (
            .O(N__11721),
            .I(\Lab_UT.scdp.prng_lfsr_3 ));
    CascadeMux I__1818 (
            .O(N__11718),
            .I(N__11715));
    InMux I__1817 (
            .O(N__11715),
            .I(N__11712));
    LocalMux I__1816 (
            .O(N__11712),
            .I(N__11709));
    Span4Mux_v I__1815 (
            .O(N__11709),
            .I(N__11706));
    Odrv4 I__1814 (
            .O(N__11706),
            .I(\Lab_UT.scdp.byteToEncrypt_3 ));
    InMux I__1813 (
            .O(N__11703),
            .I(N__11700));
    LocalMux I__1812 (
            .O(N__11700),
            .I(\Lab_UT.scdp.d2eData_3_0_3 ));
    CascadeMux I__1811 (
            .O(N__11697),
            .I(N__11694));
    InMux I__1810 (
            .O(N__11694),
            .I(N__11687));
    InMux I__1809 (
            .O(N__11693),
            .I(N__11678));
    InMux I__1808 (
            .O(N__11692),
            .I(N__11678));
    InMux I__1807 (
            .O(N__11691),
            .I(N__11678));
    InMux I__1806 (
            .O(N__11690),
            .I(N__11678));
    LocalMux I__1805 (
            .O(N__11687),
            .I(N__11673));
    LocalMux I__1804 (
            .O(N__11678),
            .I(N__11673));
    Span4Mux_v I__1803 (
            .O(N__11673),
            .I(N__11670));
    Odrv4 I__1802 (
            .O(N__11670),
            .I(\Lab_UT.scdp.N_226_i ));
    InMux I__1801 (
            .O(N__11667),
            .I(N__11664));
    LocalMux I__1800 (
            .O(N__11664),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19 ));
    CascadeMux I__1799 (
            .O(N__11661),
            .I(N__11657));
    InMux I__1798 (
            .O(N__11660),
            .I(N__11652));
    InMux I__1797 (
            .O(N__11657),
            .I(N__11648));
    InMux I__1796 (
            .O(N__11656),
            .I(N__11643));
    InMux I__1795 (
            .O(N__11655),
            .I(N__11643));
    LocalMux I__1794 (
            .O(N__11652),
            .I(N__11640));
    InMux I__1793 (
            .O(N__11651),
            .I(N__11637));
    LocalMux I__1792 (
            .O(N__11648),
            .I(\Lab_UT.scdp.d2eData_3_0_1 ));
    LocalMux I__1791 (
            .O(N__11643),
            .I(\Lab_UT.scdp.d2eData_3_0_1 ));
    Odrv12 I__1790 (
            .O(N__11640),
            .I(\Lab_UT.scdp.d2eData_3_0_1 ));
    LocalMux I__1789 (
            .O(N__11637),
            .I(\Lab_UT.scdp.d2eData_3_0_1 ));
    CascadeMux I__1788 (
            .O(N__11628),
            .I(N__11624));
    CascadeMux I__1787 (
            .O(N__11627),
            .I(N__11618));
    InMux I__1786 (
            .O(N__11624),
            .I(N__11612));
    InMux I__1785 (
            .O(N__11623),
            .I(N__11612));
    InMux I__1784 (
            .O(N__11622),
            .I(N__11607));
    InMux I__1783 (
            .O(N__11621),
            .I(N__11607));
    InMux I__1782 (
            .O(N__11618),
            .I(N__11604));
    InMux I__1781 (
            .O(N__11617),
            .I(N__11601));
    LocalMux I__1780 (
            .O(N__11612),
            .I(N__11598));
    LocalMux I__1779 (
            .O(N__11607),
            .I(N__11593));
    LocalMux I__1778 (
            .O(N__11604),
            .I(N__11593));
    LocalMux I__1777 (
            .O(N__11601),
            .I(\Lab_UT.scdp.u1.byteToDecrypt_1 ));
    Odrv4 I__1776 (
            .O(N__11598),
            .I(\Lab_UT.scdp.u1.byteToDecrypt_1 ));
    Odrv4 I__1775 (
            .O(N__11593),
            .I(\Lab_UT.scdp.u1.byteToDecrypt_1 ));
    CascadeMux I__1774 (
            .O(N__11586),
            .I(\Lab_UT.scdp.u1.N_539_cascade_ ));
    InMux I__1773 (
            .O(N__11583),
            .I(N__11580));
    LocalMux I__1772 (
            .O(N__11580),
            .I(N__11576));
    InMux I__1771 (
            .O(N__11579),
            .I(N__11571));
    Span4Mux_v I__1770 (
            .O(N__11576),
            .I(N__11568));
    InMux I__1769 (
            .O(N__11575),
            .I(N__11565));
    InMux I__1768 (
            .O(N__11574),
            .I(N__11562));
    LocalMux I__1767 (
            .O(N__11571),
            .I(\Lab_UT.scdp.N_255_i ));
    Odrv4 I__1766 (
            .O(N__11568),
            .I(\Lab_UT.scdp.N_255_i ));
    LocalMux I__1765 (
            .O(N__11565),
            .I(\Lab_UT.scdp.N_255_i ));
    LocalMux I__1764 (
            .O(N__11562),
            .I(\Lab_UT.scdp.N_255_i ));
    InMux I__1763 (
            .O(N__11553),
            .I(N__11549));
    InMux I__1762 (
            .O(N__11552),
            .I(N__11541));
    LocalMux I__1761 (
            .O(N__11549),
            .I(N__11538));
    InMux I__1760 (
            .O(N__11548),
            .I(N__11529));
    InMux I__1759 (
            .O(N__11547),
            .I(N__11529));
    InMux I__1758 (
            .O(N__11546),
            .I(N__11529));
    InMux I__1757 (
            .O(N__11545),
            .I(N__11529));
    InMux I__1756 (
            .O(N__11544),
            .I(N__11526));
    LocalMux I__1755 (
            .O(N__11541),
            .I(\Lab_UT.scdp.N_228_i ));
    Odrv4 I__1754 (
            .O(N__11538),
            .I(\Lab_UT.scdp.N_228_i ));
    LocalMux I__1753 (
            .O(N__11529),
            .I(\Lab_UT.scdp.N_228_i ));
    LocalMux I__1752 (
            .O(N__11526),
            .I(\Lab_UT.scdp.N_228_i ));
    CascadeMux I__1751 (
            .O(N__11517),
            .I(\Lab_UT.scdp.N_426_cascade_ ));
    InMux I__1750 (
            .O(N__11514),
            .I(N__11511));
    LocalMux I__1749 (
            .O(N__11511),
            .I(N__11508));
    Sp12to4 I__1748 (
            .O(N__11508),
            .I(N__11505));
    Odrv12 I__1747 (
            .O(N__11505),
            .I(\Lab_UT.scdp.q_RNI47LGA_1 ));
    InMux I__1746 (
            .O(N__11502),
            .I(N__11499));
    LocalMux I__1745 (
            .O(N__11499),
            .I(\Lab_UT.scdp.N_73 ));
    CascadeMux I__1744 (
            .O(N__11496),
            .I(\Lab_UT.scdp.N_73_cascade_ ));
    InMux I__1743 (
            .O(N__11493),
            .I(N__11490));
    LocalMux I__1742 (
            .O(N__11490),
            .I(N__11487));
    Odrv12 I__1741 (
            .O(N__11487),
            .I(\Lab_UT.scctrl.delayload ));
    InMux I__1740 (
            .O(N__11484),
            .I(N__11481));
    LocalMux I__1739 (
            .O(N__11481),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13 ));
    CascadeMux I__1738 (
            .O(N__11478),
            .I(N__11475));
    InMux I__1737 (
            .O(N__11475),
            .I(N__11472));
    LocalMux I__1736 (
            .O(N__11472),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29 ));
    InMux I__1735 (
            .O(N__11469),
            .I(N__11466));
    LocalMux I__1734 (
            .O(N__11466),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5 ));
    CascadeMux I__1733 (
            .O(N__11463),
            .I(\Lab_UT.scdp.d2eData_3_5_cascade_ ));
    InMux I__1732 (
            .O(N__11460),
            .I(N__11456));
    InMux I__1731 (
            .O(N__11459),
            .I(N__11453));
    LocalMux I__1730 (
            .O(N__11456),
            .I(N__11450));
    LocalMux I__1729 (
            .O(N__11453),
            .I(\Lab_UT.scdp.N_225_i_1 ));
    Odrv4 I__1728 (
            .O(N__11450),
            .I(\Lab_UT.scdp.N_225_i_1 ));
    InMux I__1727 (
            .O(N__11445),
            .I(N__11442));
    LocalMux I__1726 (
            .O(N__11442),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21 ));
    CascadeMux I__1725 (
            .O(N__11439),
            .I(\buart.Z_rx.N_230_cascade_ ));
    InMux I__1724 (
            .O(N__11436),
            .I(N__11433));
    LocalMux I__1723 (
            .O(N__11433),
            .I(N__11429));
    CascadeMux I__1722 (
            .O(N__11432),
            .I(N__11426));
    Span4Mux_h I__1721 (
            .O(N__11429),
            .I(N__11423));
    InMux I__1720 (
            .O(N__11426),
            .I(N__11420));
    Odrv4 I__1719 (
            .O(N__11423),
            .I(\Lab_UT.scdp.key0_7 ));
    LocalMux I__1718 (
            .O(N__11420),
            .I(\Lab_UT.scdp.key0_7 ));
    InMux I__1717 (
            .O(N__11415),
            .I(N__11412));
    LocalMux I__1716 (
            .O(N__11412),
            .I(N__11409));
    Span4Mux_v I__1715 (
            .O(N__11409),
            .I(N__11405));
    InMux I__1714 (
            .O(N__11408),
            .I(N__11402));
    Odrv4 I__1713 (
            .O(N__11405),
            .I(\Lab_UT.scdp.key0_3 ));
    LocalMux I__1712 (
            .O(N__11402),
            .I(\Lab_UT.scdp.key0_3 ));
    CascadeMux I__1711 (
            .O(N__11397),
            .I(\Lab_UT.scdp.binVal_2_cascade_ ));
    CascadeMux I__1710 (
            .O(N__11394),
            .I(\Lab_UT.scctrl.g1_0_1_cascade_ ));
    InMux I__1709 (
            .O(N__11391),
            .I(N__11388));
    LocalMux I__1708 (
            .O(N__11388),
            .I(N__11385));
    Span4Mux_v I__1707 (
            .O(N__11385),
            .I(N__11381));
    InMux I__1706 (
            .O(N__11384),
            .I(N__11378));
    Odrv4 I__1705 (
            .O(N__11381),
            .I(\Lab_UT.scdp.N_276 ));
    LocalMux I__1704 (
            .O(N__11378),
            .I(\Lab_UT.scdp.N_276 ));
    CascadeMux I__1703 (
            .O(N__11373),
            .I(N__11370));
    InMux I__1702 (
            .O(N__11370),
            .I(N__11367));
    LocalMux I__1701 (
            .O(N__11367),
            .I(N__11364));
    Span4Mux_h I__1700 (
            .O(N__11364),
            .I(N__11361));
    Odrv4 I__1699 (
            .O(N__11361),
            .I(\Lab_UT.scdp.msBitsi.N_41 ));
    InMux I__1698 (
            .O(N__11358),
            .I(N__11355));
    LocalMux I__1697 (
            .O(N__11355),
            .I(N__11352));
    Span4Mux_h I__1696 (
            .O(N__11352),
            .I(N__11349));
    Odrv4 I__1695 (
            .O(N__11349),
            .I(\ufifo.txdataDZ0Z_0 ));
    InMux I__1694 (
            .O(N__11346),
            .I(N__11343));
    LocalMux I__1693 (
            .O(N__11343),
            .I(\Lab_UT.scctrl.N_46 ));
    CascadeMux I__1692 (
            .O(N__11340),
            .I(N__11337));
    InMux I__1691 (
            .O(N__11337),
            .I(N__11334));
    LocalMux I__1690 (
            .O(N__11334),
            .I(N__11331));
    Span4Mux_s2_h I__1689 (
            .O(N__11331),
            .I(N__11328));
    Odrv4 I__1688 (
            .O(N__11328),
            .I(\buart.Z_rx.sample_i_0_a2_0 ));
    CascadeMux I__1687 (
            .O(N__11325),
            .I(N__11321));
    InMux I__1686 (
            .O(N__11324),
            .I(N__11318));
    InMux I__1685 (
            .O(N__11321),
            .I(N__11315));
    LocalMux I__1684 (
            .O(N__11318),
            .I(N__11312));
    LocalMux I__1683 (
            .O(N__11315),
            .I(\buart.Z_rx.N_230 ));
    Odrv12 I__1682 (
            .O(N__11312),
            .I(\buart.Z_rx.N_230 ));
    SRMux I__1681 (
            .O(N__11307),
            .I(N__11304));
    LocalMux I__1680 (
            .O(N__11304),
            .I(N__11298));
    CascadeMux I__1679 (
            .O(N__11303),
            .I(N__11295));
    CEMux I__1678 (
            .O(N__11302),
            .I(N__11292));
    InMux I__1677 (
            .O(N__11301),
            .I(N__11289));
    Span4Mux_v I__1676 (
            .O(N__11298),
            .I(N__11286));
    InMux I__1675 (
            .O(N__11295),
            .I(N__11283));
    LocalMux I__1674 (
            .O(N__11292),
            .I(N__11280));
    LocalMux I__1673 (
            .O(N__11289),
            .I(N__11277));
    IoSpan4Mux I__1672 (
            .O(N__11286),
            .I(N__11272));
    LocalMux I__1671 (
            .O(N__11283),
            .I(N__11272));
    Span4Mux_v I__1670 (
            .O(N__11280),
            .I(N__11269));
    Span4Mux_s1_h I__1669 (
            .O(N__11277),
            .I(N__11264));
    Span4Mux_s1_h I__1668 (
            .O(N__11272),
            .I(N__11264));
    Span4Mux_s2_h I__1667 (
            .O(N__11269),
            .I(N__11261));
    Span4Mux_h I__1666 (
            .O(N__11264),
            .I(N__11258));
    Odrv4 I__1665 (
            .O(N__11261),
            .I(\ufifo.txDataValidDZ0 ));
    Odrv4 I__1664 (
            .O(N__11258),
            .I(\ufifo.txDataValidDZ0 ));
    InMux I__1663 (
            .O(N__11253),
            .I(N__11250));
    LocalMux I__1662 (
            .O(N__11250),
            .I(N__11246));
    InMux I__1661 (
            .O(N__11249),
            .I(N__11243));
    Span4Mux_v I__1660 (
            .O(N__11246),
            .I(N__11238));
    LocalMux I__1659 (
            .O(N__11243),
            .I(N__11238));
    Odrv4 I__1658 (
            .O(N__11238),
            .I(N_233_reti));
    CascadeMux I__1657 (
            .O(N__11235),
            .I(\Lab_UT.scctrl.g1_0_1_0_cascade_ ));
    InMux I__1656 (
            .O(N__11232),
            .I(N__11225));
    InMux I__1655 (
            .O(N__11231),
            .I(N__11225));
    InMux I__1654 (
            .O(N__11230),
            .I(N__11222));
    LocalMux I__1653 (
            .O(N__11225),
            .I(\Lab_UT.sccElsBitsLd ));
    LocalMux I__1652 (
            .O(N__11222),
            .I(\Lab_UT.sccElsBitsLd ));
    CEMux I__1651 (
            .O(N__11217),
            .I(N__11213));
    CEMux I__1650 (
            .O(N__11216),
            .I(N__11210));
    LocalMux I__1649 (
            .O(N__11213),
            .I(N__11207));
    LocalMux I__1648 (
            .O(N__11210),
            .I(N__11204));
    Span4Mux_v I__1647 (
            .O(N__11207),
            .I(N__11201));
    Span4Mux_h I__1646 (
            .O(N__11204),
            .I(N__11198));
    Odrv4 I__1645 (
            .O(N__11201),
            .I(\Lab_UT.scdp.sccElsBitsLd_0 ));
    Odrv4 I__1644 (
            .O(N__11198),
            .I(\Lab_UT.scdp.sccElsBitsLd_0 ));
    InMux I__1643 (
            .O(N__11193),
            .I(N__11190));
    LocalMux I__1642 (
            .O(N__11190),
            .I(N__11187));
    Span4Mux_h I__1641 (
            .O(N__11187),
            .I(N__11184));
    Odrv4 I__1640 (
            .O(N__11184),
            .I(\Lab_UT.scdp.msBitsi.q_esr_RNI679EZ0Z_6 ));
    InMux I__1639 (
            .O(N__11181),
            .I(N__11178));
    LocalMux I__1638 (
            .O(N__11178),
            .I(N__11175));
    Odrv12 I__1637 (
            .O(N__11175),
            .I(\ufifo.txdataDZ0Z_6 ));
    InMux I__1636 (
            .O(N__11172),
            .I(N__11169));
    LocalMux I__1635 (
            .O(N__11169),
            .I(\Lab_UT.scctrl.N_534 ));
    CascadeMux I__1634 (
            .O(N__11166),
            .I(\Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0_cascade_ ));
    InMux I__1633 (
            .O(N__11163),
            .I(N__11160));
    LocalMux I__1632 (
            .O(N__11160),
            .I(\Lab_UT.scctrl.N_415_0 ));
    CascadeMux I__1631 (
            .O(N__11157),
            .I(N__11154));
    InMux I__1630 (
            .O(N__11154),
            .I(N__11151));
    LocalMux I__1629 (
            .O(N__11151),
            .I(\Lab_UT.scctrl.g1_0_0 ));
    CascadeMux I__1628 (
            .O(N__11148),
            .I(\Lab_UT.scctrl.g1_0_2_cascade_ ));
    CascadeMux I__1627 (
            .O(N__11145),
            .I(\Lab_UT.scctrl.next_state_0_0_2_cascade_ ));
    InMux I__1626 (
            .O(N__11142),
            .I(N__11139));
    LocalMux I__1625 (
            .O(N__11139),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25 ));
    InMux I__1624 (
            .O(N__11136),
            .I(N__11133));
    LocalMux I__1623 (
            .O(N__11133),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30 ));
    InMux I__1622 (
            .O(N__11130),
            .I(N__11127));
    LocalMux I__1621 (
            .O(N__11127),
            .I(N__11124));
    Odrv4 I__1620 (
            .O(N__11124),
            .I(\resetGen.N_243 ));
    InMux I__1619 (
            .O(N__11121),
            .I(N__11118));
    LocalMux I__1618 (
            .O(N__11118),
            .I(N__11115));
    Span4Mux_v I__1617 (
            .O(N__11115),
            .I(N__11112));
    Odrv4 I__1616 (
            .O(N__11112),
            .I(\buart.bu_rx_data_i_2_4 ));
    CascadeMux I__1615 (
            .O(N__11109),
            .I(N__11105));
    InMux I__1614 (
            .O(N__11108),
            .I(N__11100));
    InMux I__1613 (
            .O(N__11105),
            .I(N__11100));
    LocalMux I__1612 (
            .O(N__11100),
            .I(\Lab_UT.scdp.N_225_i_0 ));
    CascadeMux I__1611 (
            .O(N__11097),
            .I(\Lab_UT.scdp.u1.g0_0_i_a5_0_2_cascade_ ));
    InMux I__1610 (
            .O(N__11094),
            .I(N__11091));
    LocalMux I__1609 (
            .O(N__11091),
            .I(\Lab_UT.scdp.N_6 ));
    CascadeMux I__1608 (
            .O(N__11088),
            .I(\Lab_UT.scdp.u1.g0_0_i_a5_0_2_0_cascade_ ));
    InMux I__1607 (
            .O(N__11085),
            .I(N__11082));
    LocalMux I__1606 (
            .O(N__11082),
            .I(\Lab_UT.scdp.N_6_0 ));
    InMux I__1605 (
            .O(N__11079),
            .I(N__11076));
    LocalMux I__1604 (
            .O(N__11076),
            .I(N__11071));
    InMux I__1603 (
            .O(N__11075),
            .I(N__11066));
    InMux I__1602 (
            .O(N__11074),
            .I(N__11066));
    Odrv12 I__1601 (
            .O(N__11071),
            .I(\Lab_UT.scdp.d2eData_3_0_a2_0_6 ));
    LocalMux I__1600 (
            .O(N__11066),
            .I(\Lab_UT.scdp.d2eData_3_0_a2_0_6 ));
    CascadeMux I__1599 (
            .O(N__11061),
            .I(N__11056));
    CascadeMux I__1598 (
            .O(N__11060),
            .I(N__11053));
    InMux I__1597 (
            .O(N__11059),
            .I(N__11050));
    InMux I__1596 (
            .O(N__11056),
            .I(N__11045));
    InMux I__1595 (
            .O(N__11053),
            .I(N__11045));
    LocalMux I__1594 (
            .O(N__11050),
            .I(N__11042));
    LocalMux I__1593 (
            .O(N__11045),
            .I(N__11039));
    Odrv12 I__1592 (
            .O(N__11042),
            .I(\Lab_UT.scdp.prng_lfsr_14 ));
    Odrv4 I__1591 (
            .O(N__11039),
            .I(\Lab_UT.scdp.prng_lfsr_14 ));
    InMux I__1590 (
            .O(N__11034),
            .I(N__11031));
    LocalMux I__1589 (
            .O(N__11031),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17 ));
    InMux I__1588 (
            .O(N__11028),
            .I(N__11025));
    LocalMux I__1587 (
            .O(N__11025),
            .I(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22 ));
    CascadeMux I__1586 (
            .O(N__11022),
            .I(N__11019));
    InMux I__1585 (
            .O(N__11019),
            .I(N__11016));
    LocalMux I__1584 (
            .O(N__11016),
            .I(N__11013));
    Odrv4 I__1583 (
            .O(N__11013),
            .I(\Lab_UT.scdp.msBitsi.N_1919_0 ));
    InMux I__1582 (
            .O(N__11010),
            .I(N__11007));
    LocalMux I__1581 (
            .O(N__11007),
            .I(N__11004));
    Sp12to4 I__1580 (
            .O(N__11004),
            .I(N__11001));
    Odrv12 I__1579 (
            .O(N__11001),
            .I(\ufifo.txdataDZ0Z_2 ));
    CascadeMux I__1578 (
            .O(N__10998),
            .I(N__10995));
    InMux I__1577 (
            .O(N__10995),
            .I(N__10992));
    LocalMux I__1576 (
            .O(N__10992),
            .I(N__10989));
    Odrv4 I__1575 (
            .O(N__10989),
            .I(\Lab_UT.scdp.msBitsi.N_1917_0 ));
    InMux I__1574 (
            .O(N__10986),
            .I(N__10983));
    LocalMux I__1573 (
            .O(N__10983),
            .I(N__10980));
    Span4Mux_v I__1572 (
            .O(N__10980),
            .I(N__10977));
    Odrv4 I__1571 (
            .O(N__10977),
            .I(\ufifo.txdataDZ0Z_4 ));
    InMux I__1570 (
            .O(N__10974),
            .I(N__10971));
    LocalMux I__1569 (
            .O(N__10971),
            .I(\Lab_UT.scdp.N_552 ));
    CascadeMux I__1568 (
            .O(N__10968),
            .I(\Lab_UT.scdp.N_228_i_0_cascade_ ));
    InMux I__1567 (
            .O(N__10965),
            .I(N__10959));
    InMux I__1566 (
            .O(N__10964),
            .I(N__10959));
    LocalMux I__1565 (
            .O(N__10959),
            .I(N__10956));
    Odrv12 I__1564 (
            .O(N__10956),
            .I(\Lab_UT.scdp.u0.byteToDecrypt_6 ));
    InMux I__1563 (
            .O(N__10953),
            .I(N__10950));
    LocalMux I__1562 (
            .O(N__10950),
            .I(N__10947));
    Span4Mux_h I__1561 (
            .O(N__10947),
            .I(N__10944));
    Odrv4 I__1560 (
            .O(N__10944),
            .I(\Lab_UT.scdp.lfsrInst.N_234_i_0 ));
    InMux I__1559 (
            .O(N__10941),
            .I(N__10938));
    LocalMux I__1558 (
            .O(N__10938),
            .I(\Lab_UT.scdp.g0_0_i_1 ));
    CascadeMux I__1557 (
            .O(N__10935),
            .I(\Lab_UT.scdp.d2eData_3_0_1_cascade_ ));
    InMux I__1556 (
            .O(N__10932),
            .I(N__10929));
    LocalMux I__1555 (
            .O(N__10929),
            .I(\Lab_UT.scdp.msBitsi.msBitsD_1 ));
    InMux I__1554 (
            .O(N__10926),
            .I(N__10923));
    LocalMux I__1553 (
            .O(N__10923),
            .I(N__10920));
    Odrv4 I__1552 (
            .O(N__10920),
            .I(\Lab_UT.scdp.lsBitsD_1 ));
    CascadeMux I__1551 (
            .O(N__10917),
            .I(\Lab_UT.scdp.msBitsi.N_43_cascade_ ));
    InMux I__1550 (
            .O(N__10914),
            .I(N__10911));
    LocalMux I__1549 (
            .O(N__10911),
            .I(N__10908));
    Span4Mux_v I__1548 (
            .O(N__10908),
            .I(N__10905));
    Odrv4 I__1547 (
            .O(N__10905),
            .I(\ufifo.txdataDZ0Z_1 ));
    InMux I__1546 (
            .O(N__10902),
            .I(N__10899));
    LocalMux I__1545 (
            .O(N__10899),
            .I(\Lab_UT.scdp.msBitsi.msBitsD_2 ));
    InMux I__1544 (
            .O(N__10896),
            .I(N__10893));
    LocalMux I__1543 (
            .O(N__10893),
            .I(N__10890));
    Span4Mux_v I__1542 (
            .O(N__10890),
            .I(N__10887));
    Odrv4 I__1541 (
            .O(N__10887),
            .I(\Lab_UT.scdp.lsBitsD_2 ));
    InMux I__1540 (
            .O(N__10884),
            .I(N__10881));
    LocalMux I__1539 (
            .O(N__10881),
            .I(\Lab_UT.scdp.msBitsi.msBitsD_4 ));
    InMux I__1538 (
            .O(N__10878),
            .I(N__10875));
    LocalMux I__1537 (
            .O(N__10875),
            .I(N__10872));
    Odrv12 I__1536 (
            .O(N__10872),
            .I(\Lab_UT.scdp.lsBitsD_4 ));
    InMux I__1535 (
            .O(N__10869),
            .I(N__10866));
    LocalMux I__1534 (
            .O(N__10866),
            .I(N__10863));
    Span4Mux_v I__1533 (
            .O(N__10863),
            .I(N__10859));
    InMux I__1532 (
            .O(N__10862),
            .I(N__10856));
    Odrv4 I__1531 (
            .O(N__10859),
            .I(\Lab_UT.scdp.lsBitsi.lsBitsDZ0Z_5 ));
    LocalMux I__1530 (
            .O(N__10856),
            .I(\Lab_UT.scdp.lsBitsi.lsBitsDZ0Z_5 ));
    CascadeMux I__1529 (
            .O(N__10851),
            .I(\Lab_UT.scdp.N_332_i_1_cascade_ ));
    InMux I__1528 (
            .O(N__10848),
            .I(N__10845));
    LocalMux I__1527 (
            .O(N__10845),
            .I(N__10842));
    Span4Mux_v I__1526 (
            .O(N__10842),
            .I(N__10839));
    Odrv4 I__1525 (
            .O(N__10839),
            .I(\ufifo.txdataDZ0Z_5 ));
    InMux I__1524 (
            .O(N__10836),
            .I(N__10833));
    LocalMux I__1523 (
            .O(N__10833),
            .I(N__10824));
    InMux I__1522 (
            .O(N__10832),
            .I(N__10813));
    InMux I__1521 (
            .O(N__10831),
            .I(N__10813));
    InMux I__1520 (
            .O(N__10830),
            .I(N__10813));
    InMux I__1519 (
            .O(N__10829),
            .I(N__10813));
    InMux I__1518 (
            .O(N__10828),
            .I(N__10813));
    InMux I__1517 (
            .O(N__10827),
            .I(N__10810));
    Span4Mux_h I__1516 (
            .O(N__10824),
            .I(N__10807));
    LocalMux I__1515 (
            .O(N__10813),
            .I(N__10804));
    LocalMux I__1514 (
            .O(N__10810),
            .I(\Lab_UT.sccEmsBitsSl ));
    Odrv4 I__1513 (
            .O(N__10807),
            .I(\Lab_UT.sccEmsBitsSl ));
    Odrv4 I__1512 (
            .O(N__10804),
            .I(\Lab_UT.sccEmsBitsSl ));
    CascadeMux I__1511 (
            .O(N__10797),
            .I(N__10794));
    InMux I__1510 (
            .O(N__10794),
            .I(N__10791));
    LocalMux I__1509 (
            .O(N__10791),
            .I(\Lab_UT.scdp.msBitsi.msBitsD_3 ));
    InMux I__1508 (
            .O(N__10788),
            .I(N__10784));
    InMux I__1507 (
            .O(N__10787),
            .I(N__10781));
    LocalMux I__1506 (
            .O(N__10784),
            .I(N__10778));
    LocalMux I__1505 (
            .O(N__10781),
            .I(\Lab_UT.scdp.lsBitsD_3 ));
    Odrv4 I__1504 (
            .O(N__10778),
            .I(\Lab_UT.scdp.lsBitsD_3 ));
    InMux I__1503 (
            .O(N__10773),
            .I(N__10770));
    LocalMux I__1502 (
            .O(N__10770),
            .I(N__10767));
    Odrv4 I__1501 (
            .O(N__10767),
            .I(\Lab_UT.scdp.g0_0_i_1_0 ));
    InMux I__1500 (
            .O(N__10764),
            .I(N__10761));
    LocalMux I__1499 (
            .O(N__10761),
            .I(\Lab_UT.scdp.msBitsi.N_1915_0 ));
    InMux I__1498 (
            .O(N__10758),
            .I(N__10755));
    LocalMux I__1497 (
            .O(N__10755),
            .I(N__10752));
    Span4Mux_h I__1496 (
            .O(N__10752),
            .I(N__10749));
    Span4Mux_v I__1495 (
            .O(N__10749),
            .I(N__10746));
    Odrv4 I__1494 (
            .O(N__10746),
            .I(\ufifo.txdataDZ0Z_3 ));
    CascadeMux I__1493 (
            .O(N__10743),
            .I(N__10740));
    InMux I__1492 (
            .O(N__10740),
            .I(N__10737));
    LocalMux I__1491 (
            .O(N__10737),
            .I(N__10734));
    Span4Mux_h I__1490 (
            .O(N__10734),
            .I(N__10731));
    Odrv4 I__1489 (
            .O(N__10731),
            .I(\Lab_UT.scdp.byteToEncrypt_6 ));
    CascadeMux I__1488 (
            .O(N__10728),
            .I(\Lab_UT.scdp.b2a0.N_238_i_cascade_ ));
    CascadeMux I__1487 (
            .O(N__10725),
            .I(N__10719));
    CascadeMux I__1486 (
            .O(N__10724),
            .I(N__10716));
    InMux I__1485 (
            .O(N__10723),
            .I(N__10704));
    InMux I__1484 (
            .O(N__10722),
            .I(N__10704));
    InMux I__1483 (
            .O(N__10719),
            .I(N__10704));
    InMux I__1482 (
            .O(N__10716),
            .I(N__10704));
    InMux I__1481 (
            .O(N__10715),
            .I(N__10704));
    LocalMux I__1480 (
            .O(N__10704),
            .I(\Lab_UT.scdp.b2a0.N_238_i ));
    CascadeMux I__1479 (
            .O(N__10701),
            .I(N__10697));
    CascadeMux I__1478 (
            .O(N__10700),
            .I(N__10690));
    InMux I__1477 (
            .O(N__10697),
            .I(N__10685));
    InMux I__1476 (
            .O(N__10696),
            .I(N__10685));
    InMux I__1475 (
            .O(N__10695),
            .I(N__10676));
    InMux I__1474 (
            .O(N__10694),
            .I(N__10676));
    InMux I__1473 (
            .O(N__10693),
            .I(N__10676));
    InMux I__1472 (
            .O(N__10690),
            .I(N__10676));
    LocalMux I__1471 (
            .O(N__10685),
            .I(N__10671));
    LocalMux I__1470 (
            .O(N__10676),
            .I(N__10671));
    Span4Mux_h I__1469 (
            .O(N__10671),
            .I(N__10668));
    Odrv4 I__1468 (
            .O(N__10668),
            .I(\Lab_UT.scdp.b2a0.N_227_i ));
    InMux I__1467 (
            .O(N__10665),
            .I(N__10662));
    LocalMux I__1466 (
            .O(N__10662),
            .I(N__10659));
    Span4Mux_h I__1465 (
            .O(N__10659),
            .I(N__10656));
    Odrv4 I__1464 (
            .O(N__10656),
            .I(\Lab_UT.scdp.msBitsi.msBitsD_6 ));
    InMux I__1463 (
            .O(N__10653),
            .I(N__10646));
    InMux I__1462 (
            .O(N__10652),
            .I(N__10646));
    InMux I__1461 (
            .O(N__10651),
            .I(N__10643));
    LocalMux I__1460 (
            .O(N__10646),
            .I(N__10638));
    LocalMux I__1459 (
            .O(N__10643),
            .I(N__10638));
    Span4Mux_h I__1458 (
            .O(N__10638),
            .I(N__10635));
    Odrv4 I__1457 (
            .O(N__10635),
            .I(\Lab_UT.scdp.byteToEncrypt_5 ));
    InMux I__1456 (
            .O(N__10632),
            .I(N__10620));
    InMux I__1455 (
            .O(N__10631),
            .I(N__10620));
    InMux I__1454 (
            .O(N__10630),
            .I(N__10620));
    InMux I__1453 (
            .O(N__10629),
            .I(N__10620));
    LocalMux I__1452 (
            .O(N__10620),
            .I(\Lab_UT.scdp.b2a0.N_224_i ));
    InMux I__1451 (
            .O(N__10617),
            .I(N__10614));
    LocalMux I__1450 (
            .O(N__10614),
            .I(\Lab_UT.scdp.msBitsi.msBitsD_0 ));
    InMux I__1449 (
            .O(N__10611),
            .I(N__10608));
    LocalMux I__1448 (
            .O(N__10608),
            .I(N__10605));
    Odrv4 I__1447 (
            .O(N__10605),
            .I(\Lab_UT.scdp.lsBitsD_0 ));
    InMux I__1446 (
            .O(N__10602),
            .I(N__10599));
    LocalMux I__1445 (
            .O(N__10599),
            .I(N__10596));
    Span4Mux_h I__1444 (
            .O(N__10596),
            .I(N__10593));
    Odrv4 I__1443 (
            .O(N__10593),
            .I(\Lab_UT.scdp.byteToEncrypt_1 ));
    CascadeMux I__1442 (
            .O(N__10590),
            .I(N__10585));
    CascadeMux I__1441 (
            .O(N__10589),
            .I(N__10581));
    InMux I__1440 (
            .O(N__10588),
            .I(N__10572));
    InMux I__1439 (
            .O(N__10585),
            .I(N__10572));
    InMux I__1438 (
            .O(N__10584),
            .I(N__10572));
    InMux I__1437 (
            .O(N__10581),
            .I(N__10572));
    LocalMux I__1436 (
            .O(N__10572),
            .I(N__10569));
    Span4Mux_h I__1435 (
            .O(N__10569),
            .I(N__10566));
    Odrv4 I__1434 (
            .O(N__10566),
            .I(\Lab_UT.scdp.byteToEncrypt_2 ));
    CascadeMux I__1433 (
            .O(N__10563),
            .I(\Lab_UT.scdp.b2a1.N_220_i_cascade_ ));
    CascadeMux I__1432 (
            .O(N__10560),
            .I(N__10557));
    InMux I__1431 (
            .O(N__10557),
            .I(N__10545));
    InMux I__1430 (
            .O(N__10556),
            .I(N__10545));
    InMux I__1429 (
            .O(N__10555),
            .I(N__10545));
    InMux I__1428 (
            .O(N__10554),
            .I(N__10545));
    LocalMux I__1427 (
            .O(N__10545),
            .I(\Lab_UT.scdp.b2a1.N_220_i ));
    CascadeMux I__1426 (
            .O(N__10542),
            .I(\Lab_UT.scdp.N_282_cascade_ ));
    InMux I__1425 (
            .O(N__10539),
            .I(N__10533));
    InMux I__1424 (
            .O(N__10538),
            .I(N__10533));
    LocalMux I__1423 (
            .O(N__10533),
            .I(\Lab_UT.scdp.b2a1.N_293 ));
    IoInMux I__1422 (
            .O(N__10530),
            .I(N__10527));
    LocalMux I__1421 (
            .O(N__10527),
            .I(N__10523));
    InMux I__1420 (
            .O(N__10526),
            .I(N__10520));
    Span4Mux_s3_v I__1419 (
            .O(N__10523),
            .I(N__10517));
    LocalMux I__1418 (
            .O(N__10520),
            .I(N__10512));
    Span4Mux_v I__1417 (
            .O(N__10517),
            .I(N__10512));
    Odrv4 I__1416 (
            .O(N__10512),
            .I(\Lab_UT.scctrl.sccLdLFSR ));
    InMux I__1415 (
            .O(N__10509),
            .I(N__10506));
    LocalMux I__1414 (
            .O(N__10506),
            .I(\Lab_UT.scctrl.EmsLoaded ));
    CascadeMux I__1413 (
            .O(N__10503),
            .I(\Lab_UT.scctrl.EmsLoaded_cascade_ ));
    CascadeMux I__1412 (
            .O(N__10500),
            .I(\Lab_UT.sccElsBitsLd_cascade_ ));
    InMux I__1411 (
            .O(N__10497),
            .I(N__10494));
    LocalMux I__1410 (
            .O(N__10494),
            .I(\Lab_UT.scdp.lsBits_i_1_6 ));
    InMux I__1409 (
            .O(N__10491),
            .I(N__10487));
    InMux I__1408 (
            .O(N__10490),
            .I(N__10484));
    LocalMux I__1407 (
            .O(N__10487),
            .I(N__10481));
    LocalMux I__1406 (
            .O(N__10484),
            .I(\Lab_UT.scdp.lsBitsD_6 ));
    Odrv4 I__1405 (
            .O(N__10481),
            .I(\Lab_UT.scdp.lsBitsD_6 ));
    InMux I__1404 (
            .O(N__10476),
            .I(N__10472));
    InMux I__1403 (
            .O(N__10475),
            .I(N__10469));
    LocalMux I__1402 (
            .O(N__10472),
            .I(\Lab_UT.scdp.N_282 ));
    LocalMux I__1401 (
            .O(N__10469),
            .I(\Lab_UT.scdp.N_282 ));
    InMux I__1400 (
            .O(N__10464),
            .I(N__10458));
    InMux I__1399 (
            .O(N__10463),
            .I(N__10458));
    LocalMux I__1398 (
            .O(N__10458),
            .I(N__10455));
    Odrv12 I__1397 (
            .O(N__10455),
            .I(\resetGen.N_274 ));
    InMux I__1396 (
            .O(N__10452),
            .I(N__10446));
    InMux I__1395 (
            .O(N__10451),
            .I(N__10446));
    LocalMux I__1394 (
            .O(N__10446),
            .I(N__10441));
    InMux I__1393 (
            .O(N__10445),
            .I(N__10436));
    InMux I__1392 (
            .O(N__10444),
            .I(N__10436));
    Odrv12 I__1391 (
            .O(N__10441),
            .I(\resetGen.N_421 ));
    LocalMux I__1390 (
            .O(N__10436),
            .I(\resetGen.N_421 ));
    CascadeMux I__1389 (
            .O(N__10431),
            .I(N__10427));
    CascadeMux I__1388 (
            .O(N__10430),
            .I(N__10424));
    InMux I__1387 (
            .O(N__10427),
            .I(N__10419));
    InMux I__1386 (
            .O(N__10424),
            .I(N__10419));
    LocalMux I__1385 (
            .O(N__10419),
            .I(\resetGen.reset_countZ0Z_3 ));
    InMux I__1384 (
            .O(N__10416),
            .I(N__10413));
    LocalMux I__1383 (
            .O(N__10413),
            .I(N__10409));
    CascadeMux I__1382 (
            .O(N__10412),
            .I(N__10406));
    Span4Mux_v I__1381 (
            .O(N__10409),
            .I(N__10397));
    InMux I__1380 (
            .O(N__10406),
            .I(N__10394));
    InMux I__1379 (
            .O(N__10405),
            .I(N__10389));
    InMux I__1378 (
            .O(N__10404),
            .I(N__10389));
    InMux I__1377 (
            .O(N__10403),
            .I(N__10384));
    InMux I__1376 (
            .O(N__10402),
            .I(N__10384));
    InMux I__1375 (
            .O(N__10401),
            .I(N__10381));
    InMux I__1374 (
            .O(N__10400),
            .I(N__10378));
    Sp12to4 I__1373 (
            .O(N__10397),
            .I(N__10375));
    LocalMux I__1372 (
            .O(N__10394),
            .I(N__10372));
    LocalMux I__1371 (
            .O(N__10389),
            .I(N__10369));
    LocalMux I__1370 (
            .O(N__10384),
            .I(ufifo_tx_fsm_cstate_0));
    LocalMux I__1369 (
            .O(N__10381),
            .I(ufifo_tx_fsm_cstate_0));
    LocalMux I__1368 (
            .O(N__10378),
            .I(ufifo_tx_fsm_cstate_0));
    Odrv12 I__1367 (
            .O(N__10375),
            .I(ufifo_tx_fsm_cstate_0));
    Odrv4 I__1366 (
            .O(N__10372),
            .I(ufifo_tx_fsm_cstate_0));
    Odrv12 I__1365 (
            .O(N__10369),
            .I(ufifo_tx_fsm_cstate_0));
    InMux I__1364 (
            .O(N__10356),
            .I(N__10353));
    LocalMux I__1363 (
            .O(N__10353),
            .I(N__10350));
    Odrv4 I__1362 (
            .O(N__10350),
            .I(\ufifo.fifo.fifo_txdata_0 ));
    CascadeMux I__1361 (
            .O(N__10347),
            .I(N__10344));
    InMux I__1360 (
            .O(N__10344),
            .I(N__10338));
    InMux I__1359 (
            .O(N__10343),
            .I(N__10338));
    LocalMux I__1358 (
            .O(N__10338),
            .I(N__10335));
    Span4Mux_h I__1357 (
            .O(N__10335),
            .I(N__10332));
    Odrv4 I__1356 (
            .O(N__10332),
            .I(\Lab_UT.scdp.byteToEncrypt_0 ));
    InMux I__1355 (
            .O(N__10329),
            .I(\ufifo.fifo.un1_rdaddr_cry_5 ));
    CascadeMux I__1354 (
            .O(N__10326),
            .I(N__10323));
    InMux I__1353 (
            .O(N__10323),
            .I(N__10318));
    InMux I__1352 (
            .O(N__10322),
            .I(N__10315));
    InMux I__1351 (
            .O(N__10321),
            .I(N__10312));
    LocalMux I__1350 (
            .O(N__10318),
            .I(N__10307));
    LocalMux I__1349 (
            .O(N__10315),
            .I(N__10307));
    LocalMux I__1348 (
            .O(N__10312),
            .I(N__10302));
    Span4Mux_v I__1347 (
            .O(N__10307),
            .I(N__10302));
    Odrv4 I__1346 (
            .O(N__10302),
            .I(\ufifo.fifo.rdaddrZ0Z_7 ));
    InMux I__1345 (
            .O(N__10299),
            .I(\ufifo.fifo.un1_rdaddr_cry_6 ));
    InMux I__1344 (
            .O(N__10296),
            .I(bfn_4_5_0_));
    CascadeMux I__1343 (
            .O(N__10293),
            .I(N__10289));
    InMux I__1342 (
            .O(N__10292),
            .I(N__10285));
    InMux I__1341 (
            .O(N__10289),
            .I(N__10282));
    InMux I__1340 (
            .O(N__10288),
            .I(N__10279));
    LocalMux I__1339 (
            .O(N__10285),
            .I(N__10276));
    LocalMux I__1338 (
            .O(N__10282),
            .I(\ufifo.fifo.rdaddrZ0Z_8 ));
    LocalMux I__1337 (
            .O(N__10279),
            .I(\ufifo.fifo.rdaddrZ0Z_8 ));
    Odrv4 I__1336 (
            .O(N__10276),
            .I(\ufifo.fifo.rdaddrZ0Z_8 ));
    InMux I__1335 (
            .O(N__10269),
            .I(N__10264));
    InMux I__1334 (
            .O(N__10268),
            .I(N__10259));
    InMux I__1333 (
            .O(N__10267),
            .I(N__10259));
    LocalMux I__1332 (
            .O(N__10264),
            .I(N__10256));
    LocalMux I__1331 (
            .O(N__10259),
            .I(N__10253));
    Span4Mux_s3_h I__1330 (
            .O(N__10256),
            .I(N__10250));
    Odrv4 I__1329 (
            .O(N__10253),
            .I(N_251));
    Odrv4 I__1328 (
            .O(N__10250),
            .I(N_251));
    InMux I__1327 (
            .O(N__10245),
            .I(N__10242));
    LocalMux I__1326 (
            .O(N__10242),
            .I(\ufifo.fifo.fifo_txdata_1 ));
    InMux I__1325 (
            .O(N__10239),
            .I(N__10236));
    LocalMux I__1324 (
            .O(N__10236),
            .I(N__10233));
    Span4Mux_v I__1323 (
            .O(N__10233),
            .I(N__10230));
    Odrv4 I__1322 (
            .O(N__10230),
            .I(\ufifo.sb_ram512x8_inst_RNIKRN11 ));
    InMux I__1321 (
            .O(N__10227),
            .I(N__10224));
    LocalMux I__1320 (
            .O(N__10224),
            .I(N__10220));
    InMux I__1319 (
            .O(N__10223),
            .I(N__10217));
    Span4Mux_s3_h I__1318 (
            .O(N__10220),
            .I(N__10214));
    LocalMux I__1317 (
            .O(N__10217),
            .I(N__10211));
    Odrv4 I__1316 (
            .O(N__10214),
            .I(ufifo_fifo_txdata_rdy));
    Odrv4 I__1315 (
            .O(N__10211),
            .I(ufifo_fifo_txdata_rdy));
    CascadeMux I__1314 (
            .O(N__10206),
            .I(N__10202));
    InMux I__1313 (
            .O(N__10205),
            .I(N__10199));
    InMux I__1312 (
            .O(N__10202),
            .I(N__10196));
    LocalMux I__1311 (
            .O(N__10199),
            .I(N__10193));
    LocalMux I__1310 (
            .O(N__10196),
            .I(N__10190));
    Span4Mux_s3_h I__1309 (
            .O(N__10193),
            .I(N__10187));
    Odrv12 I__1308 (
            .O(N__10190),
            .I(\buart.Z_tx.N_278 ));
    Odrv4 I__1307 (
            .O(N__10187),
            .I(\buart.Z_tx.N_278 ));
    InMux I__1306 (
            .O(N__10182),
            .I(N__10170));
    InMux I__1305 (
            .O(N__10181),
            .I(N__10170));
    InMux I__1304 (
            .O(N__10180),
            .I(N__10170));
    InMux I__1303 (
            .O(N__10179),
            .I(N__10170));
    LocalMux I__1302 (
            .O(N__10170),
            .I(\resetGen.reset_countZ0Z_0 ));
    CascadeMux I__1301 (
            .O(N__10167),
            .I(N__10164));
    InMux I__1300 (
            .O(N__10164),
            .I(N__10155));
    InMux I__1299 (
            .O(N__10163),
            .I(N__10155));
    InMux I__1298 (
            .O(N__10162),
            .I(N__10155));
    LocalMux I__1297 (
            .O(N__10155),
            .I(\resetGen.reset_countZ0Z_1 ));
    InMux I__1296 (
            .O(N__10152),
            .I(N__10148));
    InMux I__1295 (
            .O(N__10151),
            .I(N__10145));
    LocalMux I__1294 (
            .O(N__10148),
            .I(\resetGen.reset_countZ0Z_2 ));
    LocalMux I__1293 (
            .O(N__10145),
            .I(\resetGen.reset_countZ0Z_2 ));
    CEMux I__1292 (
            .O(N__10140),
            .I(N__10136));
    CascadeMux I__1291 (
            .O(N__10139),
            .I(N__10131));
    LocalMux I__1290 (
            .O(N__10136),
            .I(N__10127));
    InMux I__1289 (
            .O(N__10135),
            .I(N__10124));
    InMux I__1288 (
            .O(N__10134),
            .I(N__10121));
    InMux I__1287 (
            .O(N__10131),
            .I(N__10118));
    SRMux I__1286 (
            .O(N__10130),
            .I(N__10115));
    Span4Mux_v I__1285 (
            .O(N__10127),
            .I(N__10112));
    LocalMux I__1284 (
            .O(N__10124),
            .I(N__10109));
    LocalMux I__1283 (
            .O(N__10121),
            .I(N__10104));
    LocalMux I__1282 (
            .O(N__10118),
            .I(N__10104));
    LocalMux I__1281 (
            .O(N__10115),
            .I(N__10099));
    Span4Mux_s2_h I__1280 (
            .O(N__10112),
            .I(N__10099));
    Span4Mux_h I__1279 (
            .O(N__10109),
            .I(N__10096));
    Span4Mux_h I__1278 (
            .O(N__10104),
            .I(N__10093));
    Odrv4 I__1277 (
            .O(N__10099),
            .I(\ufifo.popFifo ));
    Odrv4 I__1276 (
            .O(N__10096),
            .I(\ufifo.popFifo ));
    Odrv4 I__1275 (
            .O(N__10093),
            .I(\ufifo.popFifo ));
    CascadeMux I__1274 (
            .O(N__10086),
            .I(N__10082));
    InMux I__1273 (
            .O(N__10085),
            .I(N__10079));
    InMux I__1272 (
            .O(N__10082),
            .I(N__10076));
    LocalMux I__1271 (
            .O(N__10079),
            .I(N__10072));
    LocalMux I__1270 (
            .O(N__10076),
            .I(N__10069));
    InMux I__1269 (
            .O(N__10075),
            .I(N__10066));
    Span4Mux_s3_h I__1268 (
            .O(N__10072),
            .I(N__10063));
    Odrv4 I__1267 (
            .O(N__10069),
            .I(\ufifo.fifo.rdaddrZ0Z_0 ));
    LocalMux I__1266 (
            .O(N__10066),
            .I(\ufifo.fifo.rdaddrZ0Z_0 ));
    Odrv4 I__1265 (
            .O(N__10063),
            .I(\ufifo.fifo.rdaddrZ0Z_0 ));
    CascadeMux I__1264 (
            .O(N__10056),
            .I(N__10053));
    InMux I__1263 (
            .O(N__10053),
            .I(N__10050));
    LocalMux I__1262 (
            .O(N__10050),
            .I(N__10046));
    InMux I__1261 (
            .O(N__10049),
            .I(N__10043));
    Span4Mux_v I__1260 (
            .O(N__10046),
            .I(N__10037));
    LocalMux I__1259 (
            .O(N__10043),
            .I(N__10037));
    InMux I__1258 (
            .O(N__10042),
            .I(N__10034));
    Span4Mux_s3_h I__1257 (
            .O(N__10037),
            .I(N__10031));
    LocalMux I__1256 (
            .O(N__10034),
            .I(\ufifo.fifo.rdaddrZ0Z_1 ));
    Odrv4 I__1255 (
            .O(N__10031),
            .I(\ufifo.fifo.rdaddrZ0Z_1 ));
    InMux I__1254 (
            .O(N__10026),
            .I(\ufifo.fifo.un1_rdaddr_cry_0 ));
    CascadeMux I__1253 (
            .O(N__10023),
            .I(N__10019));
    InMux I__1252 (
            .O(N__10022),
            .I(N__10016));
    InMux I__1251 (
            .O(N__10019),
            .I(N__10013));
    LocalMux I__1250 (
            .O(N__10016),
            .I(N__10009));
    LocalMux I__1249 (
            .O(N__10013),
            .I(N__10006));
    InMux I__1248 (
            .O(N__10012),
            .I(N__10003));
    Span4Mux_s3_h I__1247 (
            .O(N__10009),
            .I(N__10000));
    Odrv4 I__1246 (
            .O(N__10006),
            .I(\ufifo.fifo.rdaddrZ0Z_2 ));
    LocalMux I__1245 (
            .O(N__10003),
            .I(\ufifo.fifo.rdaddrZ0Z_2 ));
    Odrv4 I__1244 (
            .O(N__10000),
            .I(\ufifo.fifo.rdaddrZ0Z_2 ));
    InMux I__1243 (
            .O(N__9993),
            .I(\ufifo.fifo.un1_rdaddr_cry_1 ));
    CascadeMux I__1242 (
            .O(N__9990),
            .I(N__9987));
    InMux I__1241 (
            .O(N__9987),
            .I(N__9983));
    InMux I__1240 (
            .O(N__9986),
            .I(N__9980));
    LocalMux I__1239 (
            .O(N__9983),
            .I(N__9976));
    LocalMux I__1238 (
            .O(N__9980),
            .I(N__9973));
    InMux I__1237 (
            .O(N__9979),
            .I(N__9970));
    Span4Mux_v I__1236 (
            .O(N__9976),
            .I(N__9965));
    Span4Mux_s3_h I__1235 (
            .O(N__9973),
            .I(N__9965));
    LocalMux I__1234 (
            .O(N__9970),
            .I(\ufifo.fifo.rdaddrZ0Z_3 ));
    Odrv4 I__1233 (
            .O(N__9965),
            .I(\ufifo.fifo.rdaddrZ0Z_3 ));
    InMux I__1232 (
            .O(N__9960),
            .I(\ufifo.fifo.un1_rdaddr_cry_2 ));
    CascadeMux I__1231 (
            .O(N__9957),
            .I(N__9954));
    InMux I__1230 (
            .O(N__9954),
            .I(N__9950));
    InMux I__1229 (
            .O(N__9953),
            .I(N__9947));
    LocalMux I__1228 (
            .O(N__9950),
            .I(N__9941));
    LocalMux I__1227 (
            .O(N__9947),
            .I(N__9941));
    InMux I__1226 (
            .O(N__9946),
            .I(N__9938));
    Span4Mux_s3_h I__1225 (
            .O(N__9941),
            .I(N__9935));
    LocalMux I__1224 (
            .O(N__9938),
            .I(\ufifo.fifo.rdaddrZ0Z_4 ));
    Odrv4 I__1223 (
            .O(N__9935),
            .I(\ufifo.fifo.rdaddrZ0Z_4 ));
    InMux I__1222 (
            .O(N__9930),
            .I(\ufifo.fifo.un1_rdaddr_cry_3 ));
    CascadeMux I__1221 (
            .O(N__9927),
            .I(N__9923));
    InMux I__1220 (
            .O(N__9926),
            .I(N__9920));
    InMux I__1219 (
            .O(N__9923),
            .I(N__9916));
    LocalMux I__1218 (
            .O(N__9920),
            .I(N__9913));
    InMux I__1217 (
            .O(N__9919),
            .I(N__9910));
    LocalMux I__1216 (
            .O(N__9916),
            .I(N__9905));
    Span4Mux_s3_h I__1215 (
            .O(N__9913),
            .I(N__9905));
    LocalMux I__1214 (
            .O(N__9910),
            .I(\ufifo.fifo.rdaddrZ0Z_5 ));
    Odrv4 I__1213 (
            .O(N__9905),
            .I(\ufifo.fifo.rdaddrZ0Z_5 ));
    InMux I__1212 (
            .O(N__9900),
            .I(\ufifo.fifo.un1_rdaddr_cry_4 ));
    CascadeMux I__1211 (
            .O(N__9897),
            .I(N__9894));
    InMux I__1210 (
            .O(N__9894),
            .I(N__9890));
    InMux I__1209 (
            .O(N__9893),
            .I(N__9887));
    LocalMux I__1208 (
            .O(N__9890),
            .I(N__9883));
    LocalMux I__1207 (
            .O(N__9887),
            .I(N__9880));
    InMux I__1206 (
            .O(N__9886),
            .I(N__9877));
    Span4Mux_s3_h I__1205 (
            .O(N__9883),
            .I(N__9872));
    Span4Mux_s3_h I__1204 (
            .O(N__9880),
            .I(N__9872));
    LocalMux I__1203 (
            .O(N__9877),
            .I(\ufifo.fifo.rdaddrZ0Z_6 ));
    Odrv4 I__1202 (
            .O(N__9872),
            .I(\ufifo.fifo.rdaddrZ0Z_6 ));
    InMux I__1201 (
            .O(N__9867),
            .I(N__9864));
    LocalMux I__1200 (
            .O(N__9864),
            .I(N__9861));
    IoSpan4Mux I__1199 (
            .O(N__9861),
            .I(N__9858));
    Odrv4 I__1198 (
            .O(N__9858),
            .I(uart_RXD));
    CascadeMux I__1197 (
            .O(N__9855),
            .I(N__9849));
    InMux I__1196 (
            .O(N__9854),
            .I(N__9840));
    InMux I__1195 (
            .O(N__9853),
            .I(N__9840));
    InMux I__1194 (
            .O(N__9852),
            .I(N__9840));
    InMux I__1193 (
            .O(N__9849),
            .I(N__9840));
    LocalMux I__1192 (
            .O(N__9840),
            .I(N__9837));
    Odrv4 I__1191 (
            .O(N__9837),
            .I(\Lab_UT.scdp.prng_lfsr_23 ));
    CascadeMux I__1190 (
            .O(N__9834),
            .I(\resetGen.N_421_cascade_ ));
    InMux I__1189 (
            .O(N__9831),
            .I(N__9819));
    InMux I__1188 (
            .O(N__9830),
            .I(N__9819));
    InMux I__1187 (
            .O(N__9829),
            .I(N__9819));
    InMux I__1186 (
            .O(N__9828),
            .I(N__9819));
    LocalMux I__1185 (
            .O(N__9819),
            .I(N__9816));
    Odrv4 I__1184 (
            .O(N__9816),
            .I(\buart.Z_tx.N_554 ));
    CascadeMux I__1183 (
            .O(N__9813),
            .I(\resetGen.N_267_cascade_ ));
    CascadeMux I__1182 (
            .O(N__9810),
            .I(N__9807));
    InMux I__1181 (
            .O(N__9807),
            .I(N__9804));
    LocalMux I__1180 (
            .O(N__9804),
            .I(\Lab_UT.scdp.byteToEncrypt_7 ));
    CascadeMux I__1179 (
            .O(N__9801),
            .I(N__9796));
    CascadeMux I__1178 (
            .O(N__9800),
            .I(N__9793));
    InMux I__1177 (
            .O(N__9799),
            .I(N__9783));
    InMux I__1176 (
            .O(N__9796),
            .I(N__9783));
    InMux I__1175 (
            .O(N__9793),
            .I(N__9783));
    InMux I__1174 (
            .O(N__9792),
            .I(N__9783));
    LocalMux I__1173 (
            .O(N__9783),
            .I(\Lab_UT.scdp.prng_lfsr_7 ));
    InMux I__1172 (
            .O(N__9780),
            .I(N__9768));
    InMux I__1171 (
            .O(N__9779),
            .I(N__9768));
    InMux I__1170 (
            .O(N__9778),
            .I(N__9768));
    InMux I__1169 (
            .O(N__9777),
            .I(N__9768));
    LocalMux I__1168 (
            .O(N__9768),
            .I(\Lab_UT.scdp.prng_lfsr_15 ));
    CascadeMux I__1167 (
            .O(N__9765),
            .I(\Lab_UT.scdp.lfsrInst.N_234_i_1_cascade_ ));
    InMux I__1166 (
            .O(N__9762),
            .I(N__9759));
    LocalMux I__1165 (
            .O(N__9759),
            .I(N__9756));
    Odrv4 I__1164 (
            .O(N__9756),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    InMux I__1163 (
            .O(N__9753),
            .I(N__9748));
    InMux I__1162 (
            .O(N__9752),
            .I(N__9745));
    InMux I__1161 (
            .O(N__9751),
            .I(N__9742));
    LocalMux I__1160 (
            .O(N__9748),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__1159 (
            .O(N__9745),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__1158 (
            .O(N__9742),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    InMux I__1157 (
            .O(N__9735),
            .I(N__9732));
    LocalMux I__1156 (
            .O(N__9732),
            .I(N__9729));
    Odrv4 I__1155 (
            .O(N__9729),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    InMux I__1154 (
            .O(N__9726),
            .I(N__9721));
    InMux I__1153 (
            .O(N__9725),
            .I(N__9718));
    InMux I__1152 (
            .O(N__9724),
            .I(N__9715));
    LocalMux I__1151 (
            .O(N__9721),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__1150 (
            .O(N__9718),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__1149 (
            .O(N__9715),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    InMux I__1148 (
            .O(N__9708),
            .I(N__9702));
    InMux I__1147 (
            .O(N__9707),
            .I(N__9699));
    InMux I__1146 (
            .O(N__9706),
            .I(N__9694));
    InMux I__1145 (
            .O(N__9705),
            .I(N__9694));
    LocalMux I__1144 (
            .O(N__9702),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1143 (
            .O(N__9699),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1142 (
            .O(N__9694),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__1141 (
            .O(N__9687),
            .I(N__9684));
    InMux I__1140 (
            .O(N__9684),
            .I(N__9681));
    LocalMux I__1139 (
            .O(N__9681),
            .I(N__9674));
    InMux I__1138 (
            .O(N__9680),
            .I(N__9665));
    InMux I__1137 (
            .O(N__9679),
            .I(N__9665));
    InMux I__1136 (
            .O(N__9678),
            .I(N__9665));
    InMux I__1135 (
            .O(N__9677),
            .I(N__9665));
    Odrv4 I__1134 (
            .O(N__9674),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__1133 (
            .O(N__9665),
            .I(\buart.Z_rx.ser_clk ));
    IoInMux I__1132 (
            .O(N__9660),
            .I(N__9657));
    LocalMux I__1131 (
            .O(N__9657),
            .I(N__9654));
    Span4Mux_s1_h I__1130 (
            .O(N__9654),
            .I(N__9651));
    Odrv4 I__1129 (
            .O(N__9651),
            .I(\buart.Z_rx.N_76_i ));
    InMux I__1128 (
            .O(N__9648),
            .I(N__9645));
    LocalMux I__1127 (
            .O(N__9645),
            .I(N__9642));
    Odrv4 I__1126 (
            .O(N__9642),
            .I(\ufifo.fifo.fifo_txdata_2 ));
    InMux I__1125 (
            .O(N__9639),
            .I(N__9636));
    LocalMux I__1124 (
            .O(N__9636),
            .I(N__9633));
    Odrv12 I__1123 (
            .O(N__9633),
            .I(\ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0 ));
    CascadeMux I__1122 (
            .O(N__9630),
            .I(\ufifo.sb_ram512x8_inst_RNILSN11_cascade_ ));
    InMux I__1121 (
            .O(N__9627),
            .I(N__9624));
    LocalMux I__1120 (
            .O(N__9624),
            .I(N__9621));
    Odrv12 I__1119 (
            .O(N__9621),
            .I(utb_txdata_2));
    InMux I__1118 (
            .O(N__9618),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__1117 (
            .O(N__9615),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__1116 (
            .O(N__9612),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    InMux I__1115 (
            .O(N__9609),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    CascadeMux I__1114 (
            .O(N__9606),
            .I(N__9603));
    InMux I__1113 (
            .O(N__9603),
            .I(N__9597));
    InMux I__1112 (
            .O(N__9602),
            .I(N__9597));
    LocalMux I__1111 (
            .O(N__9597),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    CascadeMux I__1110 (
            .O(N__9594),
            .I(N__9590));
    InMux I__1109 (
            .O(N__9593),
            .I(N__9585));
    InMux I__1108 (
            .O(N__9590),
            .I(N__9585));
    LocalMux I__1107 (
            .O(N__9585),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__1106 (
            .O(N__9582),
            .I(N__9578));
    InMux I__1105 (
            .O(N__9581),
            .I(N__9574));
    InMux I__1104 (
            .O(N__9578),
            .I(N__9569));
    InMux I__1103 (
            .O(N__9577),
            .I(N__9569));
    LocalMux I__1102 (
            .O(N__9574),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1101 (
            .O(N__9569),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    InMux I__1100 (
            .O(N__9564),
            .I(N__9561));
    LocalMux I__1099 (
            .O(N__9561),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3 ));
    InMux I__1098 (
            .O(N__9558),
            .I(N__9544));
    InMux I__1097 (
            .O(N__9557),
            .I(N__9544));
    InMux I__1096 (
            .O(N__9556),
            .I(N__9544));
    InMux I__1095 (
            .O(N__9555),
            .I(N__9532));
    InMux I__1094 (
            .O(N__9554),
            .I(N__9532));
    InMux I__1093 (
            .O(N__9553),
            .I(N__9532));
    InMux I__1092 (
            .O(N__9552),
            .I(N__9532));
    InMux I__1091 (
            .O(N__9551),
            .I(N__9532));
    LocalMux I__1090 (
            .O(N__9544),
            .I(N__9524));
    InMux I__1089 (
            .O(N__9543),
            .I(N__9521));
    LocalMux I__1088 (
            .O(N__9532),
            .I(N__9518));
    InMux I__1087 (
            .O(N__9531),
            .I(N__9515));
    InMux I__1086 (
            .O(N__9530),
            .I(N__9506));
    InMux I__1085 (
            .O(N__9529),
            .I(N__9506));
    InMux I__1084 (
            .O(N__9528),
            .I(N__9506));
    InMux I__1083 (
            .O(N__9527),
            .I(N__9506));
    Odrv4 I__1082 (
            .O(N__9524),
            .I(buart__tx_uart_busy_0));
    LocalMux I__1081 (
            .O(N__9521),
            .I(buart__tx_uart_busy_0));
    Odrv4 I__1080 (
            .O(N__9518),
            .I(buart__tx_uart_busy_0));
    LocalMux I__1079 (
            .O(N__9515),
            .I(buart__tx_uart_busy_0));
    LocalMux I__1078 (
            .O(N__9506),
            .I(buart__tx_uart_busy_0));
    CascadeMux I__1077 (
            .O(N__9495),
            .I(N__9492));
    InMux I__1076 (
            .O(N__9492),
            .I(N__9479));
    InMux I__1075 (
            .O(N__9491),
            .I(N__9479));
    InMux I__1074 (
            .O(N__9490),
            .I(N__9479));
    InMux I__1073 (
            .O(N__9489),
            .I(N__9479));
    InMux I__1072 (
            .O(N__9488),
            .I(N__9474));
    LocalMux I__1071 (
            .O(N__9479),
            .I(N__9471));
    InMux I__1070 (
            .O(N__9478),
            .I(N__9466));
    InMux I__1069 (
            .O(N__9477),
            .I(N__9466));
    LocalMux I__1068 (
            .O(N__9474),
            .I(\ufifo.cstate_4 ));
    Odrv4 I__1067 (
            .O(N__9471),
            .I(\ufifo.cstate_4 ));
    LocalMux I__1066 (
            .O(N__9466),
            .I(\ufifo.cstate_4 ));
    CascadeMux I__1065 (
            .O(N__9459),
            .I(\ufifo.tx_fsm.N_394_cascade_ ));
    CascadeMux I__1064 (
            .O(N__9456),
            .I(N__9453));
    InMux I__1063 (
            .O(N__9453),
            .I(N__9450));
    LocalMux I__1062 (
            .O(N__9450),
            .I(N__9447));
    Span4Mux_h I__1061 (
            .O(N__9447),
            .I(N__9442));
    InMux I__1060 (
            .O(N__9446),
            .I(N__9439));
    InMux I__1059 (
            .O(N__9445),
            .I(N__9436));
    Odrv4 I__1058 (
            .O(N__9442),
            .I(\ufifo.fifo.wraddrZ0Z_4 ));
    LocalMux I__1057 (
            .O(N__9439),
            .I(\ufifo.fifo.wraddrZ0Z_4 ));
    LocalMux I__1056 (
            .O(N__9436),
            .I(\ufifo.fifo.wraddrZ0Z_4 ));
    CascadeMux I__1055 (
            .O(N__9429),
            .I(N__9426));
    InMux I__1054 (
            .O(N__9426),
            .I(N__9423));
    LocalMux I__1053 (
            .O(N__9423),
            .I(N__9419));
    CascadeMux I__1052 (
            .O(N__9422),
            .I(N__9415));
    Span4Mux_h I__1051 (
            .O(N__9419),
            .I(N__9412));
    InMux I__1050 (
            .O(N__9418),
            .I(N__9409));
    InMux I__1049 (
            .O(N__9415),
            .I(N__9406));
    Odrv4 I__1048 (
            .O(N__9412),
            .I(\ufifo.fifo.wraddrZ0Z_5 ));
    LocalMux I__1047 (
            .O(N__9409),
            .I(\ufifo.fifo.wraddrZ0Z_5 ));
    LocalMux I__1046 (
            .O(N__9406),
            .I(\ufifo.fifo.wraddrZ0Z_5 ));
    CascadeMux I__1045 (
            .O(N__9399),
            .I(N__9396));
    InMux I__1044 (
            .O(N__9396),
            .I(N__9393));
    LocalMux I__1043 (
            .O(N__9393),
            .I(N__9390));
    Span4Mux_h I__1042 (
            .O(N__9390),
            .I(N__9385));
    InMux I__1041 (
            .O(N__9389),
            .I(N__9382));
    InMux I__1040 (
            .O(N__9388),
            .I(N__9379));
    Odrv4 I__1039 (
            .O(N__9385),
            .I(\ufifo.fifo.wraddrZ0Z_6 ));
    LocalMux I__1038 (
            .O(N__9382),
            .I(\ufifo.fifo.wraddrZ0Z_6 ));
    LocalMux I__1037 (
            .O(N__9379),
            .I(\ufifo.fifo.wraddrZ0Z_6 ));
    CascadeMux I__1036 (
            .O(N__9372),
            .I(\ufifo.fifo.un1_emptyB_NE_0_cascade_ ));
    InMux I__1035 (
            .O(N__9369),
            .I(N__9366));
    LocalMux I__1034 (
            .O(N__9366),
            .I(\ufifo.fifo.un1_emptyB_NE_3 ));
    InMux I__1033 (
            .O(N__9363),
            .I(N__9360));
    LocalMux I__1032 (
            .O(N__9360),
            .I(\ufifo.fifo.un1_emptyB_NE_2 ));
    CascadeMux I__1031 (
            .O(N__9357),
            .I(\ufifo.fifo.un1_emptyB_NE_4_cascade_ ));
    InMux I__1030 (
            .O(N__9354),
            .I(N__9351));
    LocalMux I__1029 (
            .O(N__9351),
            .I(\ufifo.fifo.un1_emptyB_NE_1 ));
    CascadeMux I__1028 (
            .O(N__9348),
            .I(\ufifo.emptyB_0_cascade_ ));
    InMux I__1027 (
            .O(N__9345),
            .I(N__9341));
    InMux I__1026 (
            .O(N__9344),
            .I(N__9338));
    LocalMux I__1025 (
            .O(N__9341),
            .I(\ufifo.tx_fsm.cstateZ0Z_5 ));
    LocalMux I__1024 (
            .O(N__9338),
            .I(\ufifo.tx_fsm.cstateZ0Z_5 ));
    CascadeMux I__1023 (
            .O(N__9333),
            .I(\ufifo.tx_fsm.N_396_cascade_ ));
    InMux I__1022 (
            .O(N__9330),
            .I(N__9322));
    InMux I__1021 (
            .O(N__9329),
            .I(N__9322));
    InMux I__1020 (
            .O(N__9328),
            .I(N__9317));
    InMux I__1019 (
            .O(N__9327),
            .I(N__9317));
    LocalMux I__1018 (
            .O(N__9322),
            .I(\ufifo.tx_fsm.N_279 ));
    LocalMux I__1017 (
            .O(N__9317),
            .I(\ufifo.tx_fsm.N_279 ));
    CascadeMux I__1016 (
            .O(N__9312),
            .I(N__9308));
    InMux I__1015 (
            .O(N__9311),
            .I(N__9303));
    InMux I__1014 (
            .O(N__9308),
            .I(N__9298));
    InMux I__1013 (
            .O(N__9307),
            .I(N__9298));
    InMux I__1012 (
            .O(N__9306),
            .I(N__9295));
    LocalMux I__1011 (
            .O(N__9303),
            .I(\ufifo.emptyB_0 ));
    LocalMux I__1010 (
            .O(N__9298),
            .I(\ufifo.emptyB_0 ));
    LocalMux I__1009 (
            .O(N__9295),
            .I(\ufifo.emptyB_0 ));
    CascadeMux I__1008 (
            .O(N__9288),
            .I(\ufifo.tx_fsm.cstate_srsts_i_0_1_1_cascade_ ));
    CascadeMux I__1007 (
            .O(N__9285),
            .I(N__9280));
    CascadeMux I__1006 (
            .O(N__9284),
            .I(N__9277));
    InMux I__1005 (
            .O(N__9283),
            .I(N__9274));
    InMux I__1004 (
            .O(N__9280),
            .I(N__9271));
    InMux I__1003 (
            .O(N__9277),
            .I(N__9268));
    LocalMux I__1002 (
            .O(N__9274),
            .I(\ufifo.tx_fsm.cstateZ0Z_1 ));
    LocalMux I__1001 (
            .O(N__9271),
            .I(\ufifo.tx_fsm.cstateZ0Z_1 ));
    LocalMux I__1000 (
            .O(N__9268),
            .I(\ufifo.tx_fsm.cstateZ0Z_1 ));
    InMux I__999 (
            .O(N__9261),
            .I(N__9258));
    LocalMux I__998 (
            .O(N__9258),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    CascadeMux I__997 (
            .O(N__9255),
            .I(utb_txdata_1_cascade_));
    InMux I__996 (
            .O(N__9252),
            .I(N__9238));
    InMux I__995 (
            .O(N__9251),
            .I(N__9231));
    InMux I__994 (
            .O(N__9250),
            .I(N__9231));
    InMux I__993 (
            .O(N__9249),
            .I(N__9231));
    InMux I__992 (
            .O(N__9248),
            .I(N__9222));
    InMux I__991 (
            .O(N__9247),
            .I(N__9222));
    InMux I__990 (
            .O(N__9246),
            .I(N__9222));
    InMux I__989 (
            .O(N__9245),
            .I(N__9222));
    InMux I__988 (
            .O(N__9244),
            .I(N__9213));
    InMux I__987 (
            .O(N__9243),
            .I(N__9213));
    InMux I__986 (
            .O(N__9242),
            .I(N__9213));
    InMux I__985 (
            .O(N__9241),
            .I(N__9213));
    LocalMux I__984 (
            .O(N__9238),
            .I(N_257));
    LocalMux I__983 (
            .O(N__9231),
            .I(N_257));
    LocalMux I__982 (
            .O(N__9222),
            .I(N_257));
    LocalMux I__981 (
            .O(N__9213),
            .I(N_257));
    InMux I__980 (
            .O(N__9204),
            .I(N__9201));
    LocalMux I__979 (
            .O(N__9201),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    CEMux I__978 (
            .O(N__9198),
            .I(N__9193));
    CEMux I__977 (
            .O(N__9197),
            .I(N__9190));
    CEMux I__976 (
            .O(N__9196),
            .I(N__9187));
    LocalMux I__975 (
            .O(N__9193),
            .I(N__9184));
    LocalMux I__974 (
            .O(N__9190),
            .I(N__9181));
    LocalMux I__973 (
            .O(N__9187),
            .I(N__9178));
    Odrv4 I__972 (
            .O(N__9184),
            .I(\buart.Z_tx.N_58 ));
    Odrv4 I__971 (
            .O(N__9181),
            .I(\buart.Z_tx.N_58 ));
    Odrv4 I__970 (
            .O(N__9178),
            .I(\buart.Z_tx.N_58 ));
    CascadeMux I__969 (
            .O(N__9171),
            .I(N__9161));
    CascadeMux I__968 (
            .O(N__9170),
            .I(N__9158));
    InMux I__967 (
            .O(N__9169),
            .I(N__9153));
    InMux I__966 (
            .O(N__9168),
            .I(N__9150));
    InMux I__965 (
            .O(N__9167),
            .I(N__9143));
    InMux I__964 (
            .O(N__9166),
            .I(N__9143));
    InMux I__963 (
            .O(N__9165),
            .I(N__9143));
    InMux I__962 (
            .O(N__9164),
            .I(N__9140));
    InMux I__961 (
            .O(N__9161),
            .I(N__9131));
    InMux I__960 (
            .O(N__9158),
            .I(N__9131));
    InMux I__959 (
            .O(N__9157),
            .I(N__9131));
    InMux I__958 (
            .O(N__9156),
            .I(N__9131));
    LocalMux I__957 (
            .O(N__9153),
            .I(ufifo_emitcrlf_fsm_cstate_0));
    LocalMux I__956 (
            .O(N__9150),
            .I(ufifo_emitcrlf_fsm_cstate_0));
    LocalMux I__955 (
            .O(N__9143),
            .I(ufifo_emitcrlf_fsm_cstate_0));
    LocalMux I__954 (
            .O(N__9140),
            .I(ufifo_emitcrlf_fsm_cstate_0));
    LocalMux I__953 (
            .O(N__9131),
            .I(ufifo_emitcrlf_fsm_cstate_0));
    CascadeMux I__952 (
            .O(N__9120),
            .I(N__9113));
    CascadeMux I__951 (
            .O(N__9119),
            .I(N__9107));
    CascadeMux I__950 (
            .O(N__9118),
            .I(N__9101));
    CascadeMux I__949 (
            .O(N__9117),
            .I(N__9098));
    InMux I__948 (
            .O(N__9116),
            .I(N__9095));
    InMux I__947 (
            .O(N__9113),
            .I(N__9082));
    InMux I__946 (
            .O(N__9112),
            .I(N__9082));
    InMux I__945 (
            .O(N__9111),
            .I(N__9082));
    InMux I__944 (
            .O(N__9110),
            .I(N__9082));
    InMux I__943 (
            .O(N__9107),
            .I(N__9082));
    InMux I__942 (
            .O(N__9106),
            .I(N__9082));
    InMux I__941 (
            .O(N__9105),
            .I(N__9073));
    InMux I__940 (
            .O(N__9104),
            .I(N__9073));
    InMux I__939 (
            .O(N__9101),
            .I(N__9073));
    InMux I__938 (
            .O(N__9098),
            .I(N__9073));
    LocalMux I__937 (
            .O(N__9095),
            .I(ufifo_emitcrlf_fsm_cstate_1));
    LocalMux I__936 (
            .O(N__9082),
            .I(ufifo_emitcrlf_fsm_cstate_1));
    LocalMux I__935 (
            .O(N__9073),
            .I(ufifo_emitcrlf_fsm_cstate_1));
    CascadeMux I__934 (
            .O(N__9066),
            .I(N__9063));
    InMux I__933 (
            .O(N__9063),
            .I(N__9060));
    LocalMux I__932 (
            .O(N__9060),
            .I(N__9057));
    Span4Mux_h I__931 (
            .O(N__9057),
            .I(N__9052));
    InMux I__930 (
            .O(N__9056),
            .I(N__9049));
    InMux I__929 (
            .O(N__9055),
            .I(N__9046));
    Odrv4 I__928 (
            .O(N__9052),
            .I(\ufifo.fifo.wraddrZ0Z_2 ));
    LocalMux I__927 (
            .O(N__9049),
            .I(\ufifo.fifo.wraddrZ0Z_2 ));
    LocalMux I__926 (
            .O(N__9046),
            .I(\ufifo.fifo.wraddrZ0Z_2 ));
    CascadeMux I__925 (
            .O(N__9039),
            .I(N__9036));
    InMux I__924 (
            .O(N__9036),
            .I(N__9033));
    LocalMux I__923 (
            .O(N__9033),
            .I(N__9029));
    CascadeMux I__922 (
            .O(N__9032),
            .I(N__9025));
    Span4Mux_h I__921 (
            .O(N__9029),
            .I(N__9022));
    InMux I__920 (
            .O(N__9028),
            .I(N__9019));
    InMux I__919 (
            .O(N__9025),
            .I(N__9016));
    Odrv4 I__918 (
            .O(N__9022),
            .I(\ufifo.fifo.wraddrZ0Z_3 ));
    LocalMux I__917 (
            .O(N__9019),
            .I(\ufifo.fifo.wraddrZ0Z_3 ));
    LocalMux I__916 (
            .O(N__9016),
            .I(\ufifo.fifo.wraddrZ0Z_3 ));
    CascadeMux I__915 (
            .O(N__9009),
            .I(N__9006));
    InMux I__914 (
            .O(N__9006),
            .I(N__9003));
    LocalMux I__913 (
            .O(N__9003),
            .I(N__8999));
    InMux I__912 (
            .O(N__9002),
            .I(N__8995));
    Span4Mux_h I__911 (
            .O(N__8999),
            .I(N__8992));
    InMux I__910 (
            .O(N__8998),
            .I(N__8989));
    LocalMux I__909 (
            .O(N__8995),
            .I(N__8986));
    Odrv4 I__908 (
            .O(N__8992),
            .I(\ufifo.fifo.wraddrZ0Z_7 ));
    LocalMux I__907 (
            .O(N__8989),
            .I(\ufifo.fifo.wraddrZ0Z_7 ));
    Odrv4 I__906 (
            .O(N__8986),
            .I(\ufifo.fifo.wraddrZ0Z_7 ));
    CascadeMux I__905 (
            .O(N__8979),
            .I(N__8975));
    CascadeMux I__904 (
            .O(N__8978),
            .I(N__8972));
    InMux I__903 (
            .O(N__8975),
            .I(N__8969));
    InMux I__902 (
            .O(N__8972),
            .I(N__8966));
    LocalMux I__901 (
            .O(N__8969),
            .I(N__8960));
    LocalMux I__900 (
            .O(N__8966),
            .I(N__8960));
    InMux I__899 (
            .O(N__8965),
            .I(N__8957));
    Span4Mux_h I__898 (
            .O(N__8960),
            .I(N__8954));
    LocalMux I__897 (
            .O(N__8957),
            .I(\ufifo.fifo.wraddrZ0Z_8 ));
    Odrv4 I__896 (
            .O(N__8954),
            .I(\ufifo.fifo.wraddrZ0Z_8 ));
    CascadeMux I__895 (
            .O(N__8949),
            .I(N__8946));
    InMux I__894 (
            .O(N__8946),
            .I(N__8943));
    LocalMux I__893 (
            .O(N__8943),
            .I(N__8940));
    Span4Mux_v I__892 (
            .O(N__8940),
            .I(N__8935));
    InMux I__891 (
            .O(N__8939),
            .I(N__8932));
    InMux I__890 (
            .O(N__8938),
            .I(N__8929));
    Odrv4 I__889 (
            .O(N__8935),
            .I(\ufifo.fifo.wraddrZ0Z_0 ));
    LocalMux I__888 (
            .O(N__8932),
            .I(\ufifo.fifo.wraddrZ0Z_0 ));
    LocalMux I__887 (
            .O(N__8929),
            .I(\ufifo.fifo.wraddrZ0Z_0 ));
    CascadeMux I__886 (
            .O(N__8922),
            .I(N__8919));
    InMux I__885 (
            .O(N__8919),
            .I(N__8916));
    LocalMux I__884 (
            .O(N__8916),
            .I(N__8912));
    CascadeMux I__883 (
            .O(N__8915),
            .I(N__8908));
    Span4Mux_v I__882 (
            .O(N__8912),
            .I(N__8905));
    InMux I__881 (
            .O(N__8911),
            .I(N__8902));
    InMux I__880 (
            .O(N__8908),
            .I(N__8899));
    Odrv4 I__879 (
            .O(N__8905),
            .I(\ufifo.fifo.wraddrZ0Z_1 ));
    LocalMux I__878 (
            .O(N__8902),
            .I(\ufifo.fifo.wraddrZ0Z_1 ));
    LocalMux I__877 (
            .O(N__8899),
            .I(\ufifo.fifo.wraddrZ0Z_1 ));
    CascadeMux I__876 (
            .O(N__8892),
            .I(\ufifo.tx_fsm.N_358_cascade_ ));
    CascadeMux I__875 (
            .O(N__8889),
            .I(\buart.Z_tx.N_373_cascade_ ));
    InMux I__874 (
            .O(N__8886),
            .I(N__8883));
    LocalMux I__873 (
            .O(N__8883),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    CascadeMux I__872 (
            .O(N__8880),
            .I(N__8877));
    InMux I__871 (
            .O(N__8877),
            .I(N__8874));
    LocalMux I__870 (
            .O(N__8874),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    CascadeMux I__869 (
            .O(N__8871),
            .I(N__8868));
    InMux I__868 (
            .O(N__8868),
            .I(N__8865));
    LocalMux I__867 (
            .O(N__8865),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    InMux I__866 (
            .O(N__8862),
            .I(N__8859));
    LocalMux I__865 (
            .O(N__8859),
            .I(\buart.Z_tx.N_375 ));
    InMux I__864 (
            .O(N__8856),
            .I(N__8853));
    LocalMux I__863 (
            .O(N__8853),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    CascadeMux I__862 (
            .O(N__8850),
            .I(\buart.Z_tx.N_215_cascade_ ));
    CascadeMux I__861 (
            .O(N__8847),
            .I(N_257_cascade_));
    CascadeMux I__860 (
            .O(N__8844),
            .I(N__8841));
    InMux I__859 (
            .O(N__8841),
            .I(N__8838));
    LocalMux I__858 (
            .O(N__8838),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    CascadeMux I__857 (
            .O(N__8835),
            .I(\ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0_cascade_ ));
    InMux I__856 (
            .O(N__8832),
            .I(\ufifo.fifo.un1_wraddr_cry_6 ));
    InMux I__855 (
            .O(N__8829),
            .I(bfn_1_7_0_));
    CascadeMux I__854 (
            .O(N__8826),
            .I(N__8823));
    InMux I__853 (
            .O(N__8823),
            .I(N__8820));
    LocalMux I__852 (
            .O(N__8820),
            .I(N__8817));
    Span4Mux_s2_h I__851 (
            .O(N__8817),
            .I(N__8814));
    Odrv4 I__850 (
            .O(N__8814),
            .I(ufifo_fifo_txdata_3));
    CascadeMux I__849 (
            .O(N__8811),
            .I(\buart.Z_tx.N_369_cascade_ ));
    CascadeMux I__848 (
            .O(N__8808),
            .I(N__8805));
    InMux I__847 (
            .O(N__8805),
            .I(N__8802));
    LocalMux I__846 (
            .O(N__8802),
            .I(N__8799));
    Span4Mux_s2_h I__845 (
            .O(N__8799),
            .I(N__8796));
    Odrv4 I__844 (
            .O(N__8796),
            .I(ufifo_fifo_txdata_4));
    CascadeMux I__843 (
            .O(N__8793),
            .I(\buart.Z_tx.N_371_cascade_ ));
    InMux I__842 (
            .O(N__8790),
            .I(N__8787));
    LocalMux I__841 (
            .O(N__8787),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__840 (
            .O(N__8784),
            .I(N__8774));
    InMux I__839 (
            .O(N__8783),
            .I(N__8774));
    InMux I__838 (
            .O(N__8782),
            .I(N__8774));
    InMux I__837 (
            .O(N__8781),
            .I(N__8771));
    LocalMux I__836 (
            .O(N__8774),
            .I(N_366));
    LocalMux I__835 (
            .O(N__8771),
            .I(N_366));
    CascadeMux I__834 (
            .O(N__8766),
            .I(N__8763));
    InMux I__833 (
            .O(N__8763),
            .I(N__8760));
    LocalMux I__832 (
            .O(N__8760),
            .I(N__8757));
    Span4Mux_s2_v I__831 (
            .O(N__8757),
            .I(N__8754));
    Odrv4 I__830 (
            .O(N__8754),
            .I(ufifo_fifo_txdata_5));
    CascadeMux I__829 (
            .O(N__8751),
            .I(\ufifo.emitcrlf_fsm.N_501_cascade_ ));
    InMux I__828 (
            .O(N__8748),
            .I(N__8745));
    LocalMux I__827 (
            .O(N__8745),
            .I(\ufifo.emitcrlf_fsm.cstate_ns_i_0_0_1 ));
    InMux I__826 (
            .O(N__8742),
            .I(\ufifo.fifo.un1_wraddr_cry_0 ));
    InMux I__825 (
            .O(N__8739),
            .I(\ufifo.fifo.un1_wraddr_cry_1 ));
    InMux I__824 (
            .O(N__8736),
            .I(\ufifo.fifo.un1_wraddr_cry_2 ));
    InMux I__823 (
            .O(N__8733),
            .I(\ufifo.fifo.un1_wraddr_cry_3 ));
    InMux I__822 (
            .O(N__8730),
            .I(\ufifo.fifo.un1_wraddr_cry_4 ));
    InMux I__821 (
            .O(N__8727),
            .I(\ufifo.fifo.un1_wraddr_cry_5 ));
    InMux I__820 (
            .O(N__8724),
            .I(N__8721));
    LocalMux I__819 (
            .O(N__8721),
            .I(N__8718));
    Span4Mux_s2_h I__818 (
            .O(N__8718),
            .I(N__8715));
    Odrv4 I__817 (
            .O(N__8715),
            .I(\ufifo.fifo.fifo_txdata_7 ));
    CascadeMux I__816 (
            .O(N__8712),
            .I(N_366_cascade_));
    CascadeMux I__815 (
            .O(N__8709),
            .I(ufifo_utb_txdata_m0_7_cascade_));
    InMux I__814 (
            .O(N__8706),
            .I(N__8703));
    LocalMux I__813 (
            .O(N__8703),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    CascadeMux I__812 (
            .O(N__8700),
            .I(\ufifo.emitcrlf_fsm.cstate_ns_i_0_2_1_cascade_ ));
    InMux I__811 (
            .O(N__8697),
            .I(N__8694));
    LocalMux I__810 (
            .O(N__8694),
            .I(\ufifo.N_323 ));
    CascadeMux I__809 (
            .O(N__8691),
            .I(\buart.Z_tx.un1_bitcount_c3_cascade_ ));
    CascadeMux I__808 (
            .O(N__8688),
            .I(N__8684));
    InMux I__807 (
            .O(N__8687),
            .I(N__8679));
    InMux I__806 (
            .O(N__8684),
            .I(N__8679));
    LocalMux I__805 (
            .O(N__8679),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    CascadeMux I__804 (
            .O(N__8676),
            .I(ufifo_utb_txdata_rdy_0_i_1_cascade_));
    CascadeMux I__803 (
            .O(N__8673),
            .I(N__8668));
    InMux I__802 (
            .O(N__8672),
            .I(N__8664));
    InMux I__801 (
            .O(N__8671),
            .I(N__8657));
    InMux I__800 (
            .O(N__8668),
            .I(N__8657));
    InMux I__799 (
            .O(N__8667),
            .I(N__8657));
    LocalMux I__798 (
            .O(N__8664),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    LocalMux I__797 (
            .O(N__8657),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    InMux I__796 (
            .O(N__8652),
            .I(N__8645));
    InMux I__795 (
            .O(N__8651),
            .I(N__8636));
    InMux I__794 (
            .O(N__8650),
            .I(N__8636));
    InMux I__793 (
            .O(N__8649),
            .I(N__8636));
    InMux I__792 (
            .O(N__8648),
            .I(N__8636));
    LocalMux I__791 (
            .O(N__8645),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__790 (
            .O(N__8636),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    InMux I__789 (
            .O(N__8631),
            .I(N__8628));
    LocalMux I__788 (
            .O(N__8628),
            .I(\buart.Z_tx.un1_bitcount_c2 ));
    InMux I__787 (
            .O(N__8625),
            .I(N__8619));
    InMux I__786 (
            .O(N__8624),
            .I(N__8619));
    LocalMux I__785 (
            .O(N__8619),
            .I(ufifo_utb_txdata_rdy_0_i_1));
    InMux I__784 (
            .O(N__8616),
            .I(N__8607));
    InMux I__783 (
            .O(N__8615),
            .I(N__8607));
    InMux I__782 (
            .O(N__8614),
            .I(N__8607));
    LocalMux I__781 (
            .O(N__8607),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__780 (
            .O(N__8604),
            .I(N__8599));
    InMux I__779 (
            .O(N__8603),
            .I(N__8591));
    InMux I__778 (
            .O(N__8602),
            .I(N__8591));
    InMux I__777 (
            .O(N__8599),
            .I(N__8582));
    InMux I__776 (
            .O(N__8598),
            .I(N__8582));
    InMux I__775 (
            .O(N__8597),
            .I(N__8582));
    InMux I__774 (
            .O(N__8596),
            .I(N__8582));
    LocalMux I__773 (
            .O(N__8591),
            .I(\buart.Z_tx.counter_RNIVE1P1_0 ));
    LocalMux I__772 (
            .O(N__8582),
            .I(\buart.Z_tx.counter_RNIVE1P1_0 ));
    CascadeMux I__771 (
            .O(N__8577),
            .I(N__8574));
    InMux I__770 (
            .O(N__8574),
            .I(N__8571));
    LocalMux I__769 (
            .O(N__8571),
            .I(N__8568));
    Span4Mux_s2_h I__768 (
            .O(N__8568),
            .I(N__8565));
    Odrv4 I__767 (
            .O(N__8565),
            .I(ufifo_fifo_txdata_6));
    IoInMux I__766 (
            .O(N__8562),
            .I(N__8559));
    LocalMux I__765 (
            .O(N__8559),
            .I(N__8556));
    IoSpan4Mux I__764 (
            .O(N__8556),
            .I(N__8553));
    IoSpan4Mux I__763 (
            .O(N__8553),
            .I(N__8550));
    Odrv4 I__762 (
            .O(N__8550),
            .I(o_serial_data_c));
    InMux I__761 (
            .O(N__8547),
            .I(N__8544));
    LocalMux I__760 (
            .O(N__8544),
            .I(\buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_6 ));
    CascadeMux I__759 (
            .O(N__8541),
            .I(N__8537));
    InMux I__758 (
            .O(N__8540),
            .I(N__8532));
    InMux I__757 (
            .O(N__8537),
            .I(N__8532));
    LocalMux I__756 (
            .O(N__8532),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    CascadeMux I__755 (
            .O(N__8529),
            .I(N__8526));
    InMux I__754 (
            .O(N__8526),
            .I(N__8523));
    LocalMux I__753 (
            .O(N__8523),
            .I(\buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_5 ));
    CascadeMux I__752 (
            .O(N__8520),
            .I(N__8517));
    InMux I__751 (
            .O(N__8517),
            .I(N__8511));
    InMux I__750 (
            .O(N__8516),
            .I(N__8511));
    LocalMux I__749 (
            .O(N__8511),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    InMux I__748 (
            .O(N__8508),
            .I(N__8504));
    InMux I__747 (
            .O(N__8507),
            .I(N__8501));
    LocalMux I__746 (
            .O(N__8504),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__745 (
            .O(N__8501),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    InMux I__744 (
            .O(N__8496),
            .I(N__8491));
    InMux I__743 (
            .O(N__8495),
            .I(N__8486));
    InMux I__742 (
            .O(N__8494),
            .I(N__8486));
    LocalMux I__741 (
            .O(N__8491),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__740 (
            .O(N__8486),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__739 (
            .O(N__8481),
            .I(N__8477));
    InMux I__738 (
            .O(N__8480),
            .I(N__8473));
    InMux I__737 (
            .O(N__8477),
            .I(N__8468));
    InMux I__736 (
            .O(N__8476),
            .I(N__8468));
    LocalMux I__735 (
            .O(N__8473),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_0 ));
    LocalMux I__734 (
            .O(N__8468),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_0 ));
    CascadeMux I__733 (
            .O(N__8463),
            .I(N__8459));
    CascadeMux I__732 (
            .O(N__8462),
            .I(N__8451));
    InMux I__731 (
            .O(N__8459),
            .I(N__8440));
    InMux I__730 (
            .O(N__8458),
            .I(N__8440));
    InMux I__729 (
            .O(N__8457),
            .I(N__8440));
    InMux I__728 (
            .O(N__8456),
            .I(N__8440));
    InMux I__727 (
            .O(N__8455),
            .I(N__8440));
    InMux I__726 (
            .O(N__8454),
            .I(N__8435));
    InMux I__725 (
            .O(N__8451),
            .I(N__8435));
    LocalMux I__724 (
            .O(N__8440),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__723 (
            .O(N__8435),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    InMux I__722 (
            .O(N__8430),
            .I(N__8421));
    InMux I__721 (
            .O(N__8429),
            .I(N__8421));
    InMux I__720 (
            .O(N__8428),
            .I(N__8421));
    LocalMux I__719 (
            .O(N__8421),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    CascadeMux I__718 (
            .O(N__8418),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_0_cascade_ ));
    CascadeMux I__717 (
            .O(N__8415),
            .I(\buart.Z_tx.counter_RNIVE1P1_0_cascade_ ));
    InMux I__716 (
            .O(N__8412),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__715 (
            .O(N__8409),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__714 (
            .O(N__8406),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__713 (
            .O(N__8403),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__712 (
            .O(N__8400),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    CascadeMux I__711 (
            .O(N__8397),
            .I(N__8394));
    InMux I__710 (
            .O(N__8394),
            .I(N__8388));
    InMux I__709 (
            .O(N__8393),
            .I(N__8388));
    LocalMux I__708 (
            .O(N__8388),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    InMux I__707 (
            .O(N__8385),
            .I(N__8382));
    LocalMux I__706 (
            .O(N__8382),
            .I(\buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_3 ));
    CascadeMux I__705 (
            .O(N__8379),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4_cascade_ ));
    InMux I__704 (
            .O(N__8376),
            .I(N__8370));
    InMux I__703 (
            .O(N__8375),
            .I(N__8370));
    LocalMux I__702 (
            .O(N__8370),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    IoInMux I__701 (
            .O(N__8367),
            .I(N__8364));
    LocalMux I__700 (
            .O(N__8364),
            .I(N__8361));
    Span12Mux_s9_v I__699 (
            .O(N__8361),
            .I(N__8358));
    Odrv12 I__698 (
            .O(N__8358),
            .I(\latticehx1k_pll_inst.clk ));
    IoInMux I__697 (
            .O(N__8355),
            .I(N__8352));
    LocalMux I__696 (
            .O(N__8352),
            .I(N__8349));
    IoSpan4Mux I__695 (
            .O(N__8349),
            .I(N__8346));
    Odrv4 I__694 (
            .O(N__8346),
            .I(clk_in_c));
    defparam IN_MUX_bfv_1_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_1_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(\ufifo.fifo.un1_wraddr_cry_7 ),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_4_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_4_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(\ufifo.fifo.un1_rdaddr_cry_7 ),
            .carryinitout(bfn_4_5_0_));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__8367),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB \resetGen.rst_1_iso_RNIU3O8  (
            .USERSIGNALTOGLOBALBUFFER(N__16451),
            .GLOBALBUFFEROUTPUT(resetGen_rst_1_iso_g));
    ICE_GB \buart.Z_rx.bitcount_es_RNIV4M42_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__9660),
            .GLOBALBUFFEROUTPUT(N_76_i_g));
    ICE_GB \Lab_UT.scctrl.state_1_ret_5_RNI  (
            .USERSIGNALTOGLOBALBUFFER(N__10530),
            .GLOBALBUFFEROUTPUT(\Lab_UT.sccLdLFSR_g ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_1_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_1_0  (
            .in0(_gnd_net_),
            .in1(N__8496),
            .in2(N__8462),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_1_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_1_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_1_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_1_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_1_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8397),
            .in3(N__8412),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__21150),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNO_0_3_LC_1_1_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_RNO_0_3_LC_1_1_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNO_0_3_LC_1_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNO_0_3_LC_1_1_2  (
            .in0(_gnd_net_),
            .in1(N__8376),
            .in2(_gnd_net_),
            .in3(N__8409),
            .lcout(\buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_1_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_1_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_1_1_3  (
            .in0(_gnd_net_),
            .in1(N__8508),
            .in2(_gnd_net_),
            .in3(N__8406),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__21150),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNO_0_5_LC_1_1_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_RNO_0_5_LC_1_1_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNO_0_5_LC_1_1_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNO_0_5_LC_1_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8520),
            .in3(N__8403),
            .lcout(\buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNO_0_6_LC_1_1_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNO_0_6_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNO_0_6_LC_1_1_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNO_0_6_LC_1_1_5  (
            .in0(_gnd_net_),
            .in1(N__8540),
            .in2(_gnd_net_),
            .in3(N__8400),
            .lcout(\buart.Z_tx.Z_baudgen.counter_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIGU38_6_LC_1_1_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIGU38_6_LC_1_1_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIGU38_6_LC_1_1_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIGU38_6_LC_1_1_6  (
            .in0(N__8516),
            .in1(N__8375),
            .in2(N__8541),
            .in3(N__8393),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(\buart.Z_tx.Z_baudgen.ser_clk_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_1_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_1_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_1_7 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_1_1_7  (
            .in0(N__8480),
            .in1(N__8385),
            .in2(N__8379),
            .in3(N__8454),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21150),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_2_0 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_2_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_2_0 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_1_2_0  (
            .in0(N__8458),
            .in1(N__8547),
            .in2(N__8481),
            .in3(N__8430),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_2_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_2_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_2_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_1_2_1  (
            .in0(N__8429),
            .in1(N__8476),
            .in2(N__8529),
            .in3(N__8457),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_2_2 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_2_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_2_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_1_2_2  (
            .in0(N__8456),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_2_4 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_2_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_2_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_1_2_4  (
            .in0(N__8495),
            .in1(_gnd_net_),
            .in2(N__8463),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21149),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5S14_1_LC_1_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5S14_1_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5S14_1_LC_1_2_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5S14_1_LC_1_2_5  (
            .in0(_gnd_net_),
            .in1(N__8507),
            .in2(_gnd_net_),
            .in3(N__8494),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_0 ),
            .ltout(\buart.Z_tx.Z_baudgen.ser_clk_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_0_LC_1_2_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_0_LC_1_2_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_0_LC_1_2_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIVE1P1_0_LC_1_2_6  (
            .in0(N__8455),
            .in1(N__8428),
            .in2(N__8418),
            .in3(N__9543),
            .lcout(\buart.Z_tx.counter_RNIVE1P1_0 ),
            .ltout(\buart.Z_tx.counter_RNIVE1P1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_1_2_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_1_2_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_1_2_7 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_1_2_7  (
            .in0(_gnd_net_),
            .in1(N__8672),
            .in2(N__8415),
            .in3(N__8652),
            .lcout(\buart.Z_tx.un1_bitcount_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_1_3_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_1_3_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_tx.bitcount_RNIQOQA1_3_LC_1_3_0  (
            .in0(N__8614),
            .in1(N__8667),
            .in2(N__8688),
            .in3(N__8648),
            .lcout(buart__tx_uart_busy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_1_3_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_1_3_1 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_1_3_1  (
            .in0(N__8649),
            .in1(N__8596),
            .in2(N__8673),
            .in3(N__8615),
            .lcout(),
            .ltout(\buart.Z_tx.un1_bitcount_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_3_LC_1_3_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_1_3_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_1_3_2 .LUT_INIT=16'b1111111110010110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_1_3_2  (
            .in0(N__8687),
            .in1(N__8603),
            .in2(N__8691),
            .in3(N__8625),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21148),
            .ce(),
            .sr(N__20833));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIPKRF7_0_LC_1_3_3 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIPKRF7_0_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIPKRF7_0_LC_1_3_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIPKRF7_0_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(N__12320),
            .in2(_gnd_net_),
            .in3(N__9249),
            .lcout(ufifo_utb_txdata_rdy_0_i_1),
            .ltout(ufifo_utb_txdata_rdy_0_i_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_1_LC_1_3_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_1_3_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_1_3_4 .LUT_INIT=16'b1111110011110110;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_1_3_4  (
            .in0(N__8598),
            .in1(N__8671),
            .in2(N__8676),
            .in3(N__8650),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21148),
            .ce(),
            .sr(N__20833));
    defparam \buart.Z_tx.bitcount_0_LC_1_3_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_1_3_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_1_3_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_1_3_5  (
            .in0(N__8651),
            .in1(N__8597),
            .in2(_gnd_net_),
            .in3(N__9251),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21148),
            .ce(),
            .sr(N__20833));
    defparam \buart.Z_tx.bitcount_2_LC_1_3_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_1_3_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_1_3_6 .LUT_INIT=16'b0000000010010110;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_1_3_6  (
            .in0(N__8616),
            .in1(N__8631),
            .in2(N__8604),
            .in3(N__8624),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21148),
            .ce(),
            .sr(N__20833));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIO3T89_0_LC_1_3_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIO3T89_0_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIO3T89_0_LC_1_3_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIO3T89_0_LC_1_3_7  (
            .in0(N__8602),
            .in1(N__12321),
            .in2(_gnd_net_),
            .in3(N__9250),
            .lcout(\buart.Z_tx.N_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_RNO_0_7_LC_1_4_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_RNO_0_7_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.shifter_RNO_0_7_LC_1_4_0 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \buart.Z_tx.shifter_RNO_0_7_LC_1_4_0  (
            .in0(N__8781),
            .in1(N__14935),
            .in2(N__8577),
            .in3(N__9241),
            .lcout(\buart.Z_tx.N_375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.uart_tx_LC_1_4_1 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_1_4_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_1_4_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \buart.Z_tx.uart_tx_LC_1_4_1  (
            .in0(N__9244),
            .in1(N__8706),
            .in2(_gnd_net_),
            .in3(N__12315),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21146),
            .ce(N__9196),
            .sr(N__20831));
    defparam \ufifo.tx_fsm.cstate_RNI57IK1_0_LC_1_4_2 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNI57IK1_0_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNI57IK1_0_LC_1_4_2 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \ufifo.tx_fsm.cstate_RNI57IK1_0_LC_1_4_2  (
            .in0(N__9168),
            .in1(N__9116),
            .in2(N__10412),
            .in3(N__9531),
            .lcout(N_366),
            .ltout(N_366_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIEQME2_LC_1_4_3 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIEQME2_LC_1_4_3 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIEQME2_LC_1_4_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNIEQME2_LC_1_4_3  (
            .in0(_gnd_net_),
            .in1(N__8724),
            .in2(N__8712),
            .in3(N__14529),
            .lcout(),
            .ltout(ufifo_utb_txdata_m0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_8_LC_1_4_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_1_4_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_1_4_4 .LUT_INIT=16'b0101000001010101;
    LogicCell40 \buart.Z_tx.shifter_8_LC_1_4_4  (
            .in0(N__12314),
            .in1(_gnd_net_),
            .in2(N__8709),
            .in3(N__9243),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21146),
            .ce(N__9196),
            .sr(N__20831));
    defparam \buart.Z_tx.shifter_0_LC_1_4_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_1_4_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_1_4_5 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \buart.Z_tx.shifter_0_LC_1_4_5  (
            .in0(N__9242),
            .in1(_gnd_net_),
            .in2(N__8844),
            .in3(N__12313),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21146),
            .ce(N__9196),
            .sr(N__20831));
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_0_1_LC_1_5_0 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_0_1_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_0_1_LC_1_5_0 .LUT_INIT=16'b1111111101100100;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNO_0_1_LC_1_5_0  (
            .in0(N__9554),
            .in1(N__9111),
            .in2(N__9171),
            .in3(N__8748),
            .lcout(),
            .ltout(\ufifo.emitcrlf_fsm.cstate_ns_i_0_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_1_LC_1_5_1 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_1_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \ufifo.emitcrlf_fsm.cstate_1_LC_1_5_1 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_1_LC_1_5_1  (
            .in0(N__9112),
            .in1(N__8697),
            .in2(N__8700),
            .in3(N__15449),
            .lcout(ufifo_emitcrlf_fsm_cstate_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21144),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNI7ELR5_4_LC_1_5_2 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNI7ELR5_4_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNI7ELR5_4_LC_1_5_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \ufifo.tx_fsm.cstate_RNI7ELR5_4_LC_1_5_2  (
            .in0(N__9553),
            .in1(N__9478),
            .in2(_gnd_net_),
            .in3(N__9306),
            .lcout(\ufifo.N_323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_0_LC_1_5_3 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_0_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \ufifo.emitcrlf_fsm.cstate_0_LC_1_5_3 .LUT_INIT=16'b0110101000000000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_0_LC_1_5_3  (
            .in0(N__9169),
            .in1(N__9555),
            .in2(N__9120),
            .in3(N__15448),
            .lcout(ufifo_emitcrlf_fsm_cstate_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21144),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_srsts_i_i_o2_2_LC_1_5_4 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_srsts_i_i_o2_2_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_srsts_i_i_o2_2_LC_1_5_4 .LUT_INIT=16'b0111111101111111;
    LogicCell40 \ufifo.tx_fsm.cstate_srsts_i_i_o2_2_LC_1_5_4  (
            .in0(N__9552),
            .in1(N__9110),
            .in2(N__9170),
            .in3(_gnd_net_),
            .lcout(\ufifo.tx_fsm.N_279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_0_LC_1_5_5 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_0_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_0_LC_1_5_5 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_0_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(N__9551),
            .in2(N__9119),
            .in3(N__9156),
            .lcout(N_368),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_2_1_LC_1_5_6 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_2_1_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_2_1_LC_1_5_6 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNO_2_1_LC_1_5_6  (
            .in0(N__9157),
            .in1(N__9106),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\ufifo.emitcrlf_fsm.N_501_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_1_1_LC_1_5_7 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_1_1_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNO_1_1_LC_1_5_7 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNO_1_1_LC_1_5_7  (
            .in0(N__9477),
            .in1(N__10401),
            .in2(N__8751),
            .in3(N__23208),
            .lcout(\ufifo.emitcrlf_fsm.cstate_ns_i_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_0_LC_1_6_0 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_0_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_0_LC_1_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_0_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__8939),
            .in2(N__11303),
            .in3(N__11301),
            .lcout(\ufifo.fifo.wraddrZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\ufifo.fifo.un1_wraddr_cry_0 ),
            .clk(N__21140),
            .ce(),
            .sr(N__20808));
    defparam \ufifo.fifo.wraddr_1_LC_1_6_1 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_1_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_1_LC_1_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_1_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__8911),
            .in2(_gnd_net_),
            .in3(N__8742),
            .lcout(\ufifo.fifo.wraddrZ0Z_1 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_0 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_1 ),
            .clk(N__21140),
            .ce(),
            .sr(N__20808));
    defparam \ufifo.fifo.wraddr_2_LC_1_6_2 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_2_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_2_LC_1_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_2_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__9056),
            .in2(_gnd_net_),
            .in3(N__8739),
            .lcout(\ufifo.fifo.wraddrZ0Z_2 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_1 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_2 ),
            .clk(N__21140),
            .ce(),
            .sr(N__20808));
    defparam \ufifo.fifo.wraddr_3_LC_1_6_3 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_3_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_3_LC_1_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_3_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(N__9028),
            .in2(_gnd_net_),
            .in3(N__8736),
            .lcout(\ufifo.fifo.wraddrZ0Z_3 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_2 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_3 ),
            .clk(N__21140),
            .ce(),
            .sr(N__20808));
    defparam \ufifo.fifo.wraddr_4_LC_1_6_4 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_4_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_4_LC_1_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_4_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(N__9446),
            .in2(_gnd_net_),
            .in3(N__8733),
            .lcout(\ufifo.fifo.wraddrZ0Z_4 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_3 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_4 ),
            .clk(N__21140),
            .ce(),
            .sr(N__20808));
    defparam \ufifo.fifo.wraddr_5_LC_1_6_5 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_5_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_5_LC_1_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_5_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(N__9418),
            .in2(_gnd_net_),
            .in3(N__8730),
            .lcout(\ufifo.fifo.wraddrZ0Z_5 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_4 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_5 ),
            .clk(N__21140),
            .ce(),
            .sr(N__20808));
    defparam \ufifo.fifo.wraddr_6_LC_1_6_6 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_6_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_6_LC_1_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_6_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(N__9389),
            .in2(_gnd_net_),
            .in3(N__8727),
            .lcout(\ufifo.fifo.wraddrZ0Z_6 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_5 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_6 ),
            .clk(N__21140),
            .ce(),
            .sr(N__20808));
    defparam \ufifo.fifo.wraddr_7_LC_1_6_7 .C_ON=1'b1;
    defparam \ufifo.fifo.wraddr_7_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_7_LC_1_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.wraddr_7_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(N__8998),
            .in2(_gnd_net_),
            .in3(N__8832),
            .lcout(\ufifo.fifo.wraddrZ0Z_7 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_wraddr_cry_6 ),
            .carryout(\ufifo.fifo.un1_wraddr_cry_7 ),
            .clk(N__21140),
            .ce(),
            .sr(N__20808));
    defparam \ufifo.fifo.wraddr_8_LC_1_7_0 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_8_LC_1_7_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.wraddr_8_LC_1_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ufifo.fifo.wraddr_8_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__8965),
            .in2(_gnd_net_),
            .in3(N__8829),
            .lcout(\ufifo.fifo.wraddrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21132),
            .ce(),
            .sr(N__20807));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_1_9_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_1_9_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_1_9_6  (
            .in0(N__9705),
            .in1(N__9724),
            .in2(_gnd_net_),
            .in3(N__9564),
            .lcout(\buart.Z_rx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_1_9_7 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_1_9_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_1_9_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_1_9_7  (
            .in0(N__9581),
            .in1(N__17703),
            .in2(_gnd_net_),
            .in3(N__9706),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21121),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.EmsBitsSl_LC_1_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.EmsBitsSl_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.EmsBitsSl_LC_1_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.scctrl.EmsBitsSl_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10827),
            .lcout(\Lab_UT.sccEmsBitsSl ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21108),
            .ce(),
            .sr(N__20810));
    defparam \buart.Z_tx.shifter_RNO_0_4_LC_2_3_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_RNO_0_4_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.shifter_RNO_0_4_LC_2_3_0 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \buart.Z_tx.shifter_RNO_0_4_LC_2_3_0  (
            .in0(N__8782),
            .in1(N__13551),
            .in2(N__8826),
            .in3(N__9245),
            .lcout(),
            .ltout(\buart.Z_tx.N_369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_4_LC_2_3_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_2_3_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_2_3_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \buart.Z_tx.shifter_4_LC_2_3_1  (
            .in0(N__12322),
            .in1(N__8790),
            .in2(N__8811),
            .in3(N__9828),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__9197),
            .sr(N__20838));
    defparam \buart.Z_tx.shifter_RNO_0_5_LC_2_3_2 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_RNO_0_5_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.shifter_RNO_0_5_LC_2_3_2 .LUT_INIT=16'b0000100001001100;
    LogicCell40 \buart.Z_tx.shifter_RNO_0_5_LC_2_3_2  (
            .in0(N__8783),
            .in1(N__9246),
            .in2(N__8808),
            .in3(N__15127),
            .lcout(),
            .ltout(\buart.Z_tx.N_371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_5_LC_2_3_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_2_3_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_2_3_3 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \buart.Z_tx.shifter_5_LC_2_3_3  (
            .in0(N__12323),
            .in1(N__8886),
            .in2(N__8793),
            .in3(N__9829),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__9197),
            .sr(N__20838));
    defparam \buart.Z_tx.shifter_RNO_0_6_LC_2_3_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_RNO_0_6_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.shifter_RNO_0_6_LC_2_3_4 .LUT_INIT=16'b0000100001001100;
    LogicCell40 \buart.Z_tx.shifter_RNO_0_6_LC_2_3_4  (
            .in0(N__8784),
            .in1(N__9247),
            .in2(N__8766),
            .in3(N__18808),
            .lcout(),
            .ltout(\buart.Z_tx.N_373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_6_LC_2_3_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_2_3_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_2_3_5 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \buart.Z_tx.shifter_6_LC_2_3_5  (
            .in0(N__12324),
            .in1(N__8856),
            .in2(N__8889),
            .in3(N__9830),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__9197),
            .sr(N__20838));
    defparam \buart.Z_tx.shifter_3_LC_2_3_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_2_3_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_2_3_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \buart.Z_tx.shifter_3_LC_2_3_6  (
            .in0(N__9627),
            .in1(N__12326),
            .in2(N__8880),
            .in3(N__9248),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__9197),
            .sr(N__20838));
    defparam \buart.Z_tx.shifter_7_LC_2_3_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_2_3_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_2_3_7 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \buart.Z_tx.shifter_7_LC_2_3_7  (
            .in0(N__12325),
            .in1(N__9831),
            .in2(N__8871),
            .in3(N__8862),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21147),
            .ce(N__9197),
            .sr(N__20838));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2_0_LC_2_4_0 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2_0_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2_0_LC_2_4_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2_0_LC_2_4_0  (
            .in0(N__9529),
            .in1(N__9104),
            .in2(_gnd_net_),
            .in3(N__9165),
            .lcout(\ufifo.emitcrlf_fsm.cstate_RNIJLRB1_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIF2CB3_3_LC_2_4_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIF2CB3_3_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIF2CB3_3_LC_2_4_1 .LUT_INIT=16'b0100100011111111;
    LogicCell40 \buart.Z_tx.bitcount_RNIF2CB3_3_LC_2_4_1  (
            .in0(N__9166),
            .in1(N__9527),
            .in2(N__9117),
            .in3(N__14383),
            .lcout(),
            .ltout(\buart.Z_tx.N_215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNI6VV36_3_LC_2_4_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNI6VV36_3_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNI6VV36_3_LC_2_4_2 .LUT_INIT=16'b1111001110110011;
    LogicCell40 \buart.Z_tx.bitcount_RNI6VV36_3_LC_2_4_2  (
            .in0(N__11121),
            .in1(N__10205),
            .in2(N__8850),
            .in3(N__10269),
            .lcout(N_257),
            .ltout(N_257_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_2_4_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_2_4_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_2_4_3 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \buart.Z_tx.shifter_1_LC_2_4_3  (
            .in0(N__9204),
            .in1(N__12255),
            .in2(N__8847),
            .in3(N__12311),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21145),
            .ce(N__9198),
            .sr(N__20835));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_LC_2_4_4 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_LC_2_4_4 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_0_LC_2_4_4  (
            .in0(N__9530),
            .in1(N__9105),
            .in2(_gnd_net_),
            .in3(N__9167),
            .lcout(),
            .ltout(\ufifo.emitcrlf_fsm.cstate_RNIJLRB1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIQ6FP3_0_LC_2_4_5 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIQ6FP3_0_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIQ6FP3_0_LC_2_4_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIQ6FP3_0_LC_2_4_5  (
            .in0(_gnd_net_),
            .in1(N__10239),
            .in2(N__8835),
            .in3(N__12310),
            .lcout(),
            .ltout(utb_txdata_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_2_LC_2_4_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_2_4_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_2_4_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \buart.Z_tx.shifter_2_LC_2_4_6  (
            .in0(N__12312),
            .in1(N__9261),
            .in2(N__9255),
            .in3(N__9252),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21145),
            .ce(N__9198),
            .sr(N__20835));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1_0_LC_2_4_7 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1_0_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1_0_LC_2_4_7 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1_0_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(N__9164),
            .in2(N__9118),
            .in3(N__9528),
            .lcout(\ufifo.emitcrlf_fsm.cstate_RNIJLRB1_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_RNIOP7U_2_LC_2_5_0 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNIOP7U_2_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNIOP7U_2_LC_2_5_0 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \ufifo.fifo.wraddr_RNIOP7U_2_LC_2_5_0  (
            .in0(N__9055),
            .in1(N__9986),
            .in2(N__9032),
            .in3(N__10022),
            .lcout(\ufifo.fifo.un1_emptyB_NE_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_RNICE8U_8_LC_2_5_1 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNICE8U_8_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNICE8U_8_LC_2_5_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \ufifo.fifo.wraddr_RNICE8U_8_LC_2_5_1  (
            .in0(N__9002),
            .in1(N__10292),
            .in2(N__8978),
            .in3(N__10322),
            .lcout(\ufifo.fifo.un1_emptyB_NE_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_RNIGH7U_0_LC_2_5_2 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNIGH7U_0_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNIGH7U_0_LC_2_5_2 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \ufifo.fifo.wraddr_RNIGH7U_0_LC_2_5_2  (
            .in0(N__8938),
            .in1(N__10049),
            .in2(N__8915),
            .in3(N__10085),
            .lcout(\ufifo.fifo.un1_emptyB_NE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNO_0_2_LC_2_5_3 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNO_0_2_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNO_0_2_LC_2_5_3 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \ufifo.tx_fsm.cstate_RNO_0_2_LC_2_5_3  (
            .in0(N__9490),
            .in1(N__9307),
            .in2(N__9284),
            .in3(N__9556),
            .lcout(),
            .ltout(\ufifo.tx_fsm.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_2_LC_2_5_4 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_2_LC_2_5_4 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_2_LC_2_5_4 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \ufifo.tx_fsm.cstate_2_LC_2_5_4  (
            .in0(N__20176),
            .in1(N__9491),
            .in2(N__8892),
            .in3(N__9329),
            .lcout(\ufifo.popFifo ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_4_LC_2_5_5 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_4_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_4_LC_2_5_5 .LUT_INIT=16'b0010001000110010;
    LogicCell40 \ufifo.tx_fsm.cstate_4_LC_2_5_5  (
            .in0(N__10227),
            .in1(N__20177),
            .in2(N__9495),
            .in3(N__9558),
            .lcout(\ufifo.cstate_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNO_0_5_LC_2_5_6 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNO_0_5_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNO_0_5_LC_2_5_6 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \ufifo.tx_fsm.cstate_RNO_0_5_LC_2_5_6  (
            .in0(N__9557),
            .in1(N__9344),
            .in2(N__9312),
            .in3(N__9489),
            .lcout(),
            .ltout(\ufifo.tx_fsm.N_394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_5_LC_2_5_7 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_5_LC_2_5_7 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_5_LC_2_5_7 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \ufifo.tx_fsm.cstate_5_LC_2_5_7  (
            .in0(N__9330),
            .in1(N__9488),
            .in2(N__9459),
            .in3(N__20178),
            .lcout(\ufifo.tx_fsm.cstateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21141),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_RNI028U_4_LC_2_6_0 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNI028U_4_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNI028U_4_LC_2_6_0 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \ufifo.fifo.wraddr_RNI028U_4_LC_2_6_0  (
            .in0(N__9445),
            .in1(N__9926),
            .in2(N__9422),
            .in3(N__9953),
            .lcout(),
            .ltout(\ufifo.fifo.un1_emptyB_NE_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_RNI36CD1_6_LC_2_6_1 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNI36CD1_6_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNI36CD1_6_LC_2_6_1 .LUT_INIT=16'b1100000000110000;
    LogicCell40 \ufifo.fifo.wraddr_RNI36CD1_6_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__9388),
            .in2(N__9372),
            .in3(N__9893),
            .lcout(),
            .ltout(\ufifo.fifo.un1_emptyB_NE_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.wraddr_RNINV384_0_LC_2_6_2 .C_ON=1'b0;
    defparam \ufifo.fifo.wraddr_RNINV384_0_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.wraddr_RNINV384_0_LC_2_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ufifo.fifo.wraddr_RNINV384_0_LC_2_6_2  (
            .in0(N__9369),
            .in1(N__9363),
            .in2(N__9357),
            .in3(N__9354),
            .lcout(\ufifo.emptyB_0 ),
            .ltout(\ufifo.emptyB_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNO_0_0_LC_2_6_3 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNO_0_0_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNO_0_0_LC_2_6_3 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \ufifo.tx_fsm.cstate_RNO_0_0_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(N__10402),
            .in2(N__9348),
            .in3(N__23210),
            .lcout(),
            .ltout(\ufifo.tx_fsm.N_396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstateZ0Z_0_LC_2_6_4 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstateZ0Z_0_LC_2_6_4 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstateZ0Z_0_LC_2_6_4 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \ufifo.tx_fsm.cstateZ0Z_0_LC_2_6_4  (
            .in0(N__20175),
            .in1(N__9345),
            .in2(N__9333),
            .in3(N__9328),
            .lcout(ufifo_tx_fsm_cstate_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21133),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_RNO_0_1_LC_2_6_5 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_RNO_0_1_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \ufifo.tx_fsm.cstate_RNO_0_1_LC_2_6_5 .LUT_INIT=16'b0001000000011100;
    LogicCell40 \ufifo.tx_fsm.cstate_RNO_0_1_LC_2_6_5  (
            .in0(N__9327),
            .in1(N__10403),
            .in2(N__9285),
            .in3(N__23211),
            .lcout(),
            .ltout(\ufifo.tx_fsm.cstate_srsts_i_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_1_LC_2_6_6 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_1_LC_2_6_6 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_1_LC_2_6_6 .LUT_INIT=16'b0001101000000000;
    LogicCell40 \ufifo.tx_fsm.cstate_1_LC_2_6_6  (
            .in0(N__9283),
            .in1(N__9311),
            .in2(N__9288),
            .in3(N__15459),
            .lcout(\ufifo.tx_fsm.cstateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21133),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNILSN11_LC_2_7_1 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNILSN11_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNILSN11_LC_2_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNILSN11_LC_2_7_1  (
            .in0(N__9648),
            .in1(N__10400),
            .in2(_gnd_net_),
            .in3(N__13032),
            .lcout(),
            .ltout(\ufifo.sb_ram512x8_inst_RNILSN11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIR7FP3_0_LC_2_7_2 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIR7FP3_0_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIR7FP3_0_LC_2_7_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIR7FP3_0_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__9639),
            .in2(N__9630),
            .in3(N__12316),
            .lcout(utb_txdata_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_9_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__9707),
            .in2(N__9582),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_9_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__9725),
            .in2(_gnd_net_),
            .in3(N__9618),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_2_9_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_2_9_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_2_9_2  (
            .in0(N__17702),
            .in1(_gnd_net_),
            .in2(N__9606),
            .in3(N__9615),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__21116),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_9_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__9752),
            .in2(_gnd_net_),
            .in3(N__9612),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_2_9_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_2_9_4 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_2_9_4  (
            .in0(N__17701),
            .in1(N__9593),
            .in2(N__9687),
            .in3(N__9609),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21116),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_9_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_9_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_9_5  (
            .in0(N__9751),
            .in1(N__9602),
            .in2(N__9594),
            .in3(N__9577),
            .lcout(\buart.Z_rx.Z_baudgen.ser_clk_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_2_10_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_2_10_2 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_2_10_2  (
            .in0(N__9680),
            .in1(N__9762),
            .in2(N__17700),
            .in3(N__9753),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_10_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_10_4 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_2_10_4  (
            .in0(N__9679),
            .in1(N__9735),
            .in2(N__17699),
            .in3(N__9726),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_2_10_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_2_10_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(N__9708),
            .in2(_gnd_net_),
            .in3(N__17685),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21109),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIELQA6_0_LC_2_10_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIELQA6_0_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIELQA6_0_LC_2_10_6 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIELQA6_0_LC_2_10_6  (
            .in0(N__9678),
            .in1(N__17793),
            .in2(N__17698),
            .in3(N__14366),
            .lcout(\buart.Z_rx.N_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_10_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_10_7 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_10_7  (
            .in0(N__11324),
            .in1(N__9677),
            .in2(N__11340),
            .in3(N__13869),
            .lcout(\buart.Z_rx.N_76_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u2.q_esr_0_LC_2_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_0_LC_2_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_0_LC_2_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_0_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16580),
            .lcout(\Lab_UT.scdp.byteToEncrypt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21100),
            .ce(N__13905),
            .sr(N__20811));
    defparam \Lab_UT.scdp.u2.q_esr_1_LC_2_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_1_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_1_LC_2_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_1_LC_2_11_1  (
            .in0(N__17205),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scdp.byteToEncrypt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21100),
            .ce(N__13905),
            .sr(N__20811));
    defparam \Lab_UT.scdp.u2.q_esr_2_LC_2_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_2_LC_2_11_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_2_LC_2_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_2_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13033),
            .lcout(\Lab_UT.scdp.byteToEncrypt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21100),
            .ce(N__13905),
            .sr(N__20811));
    defparam \Lab_UT.scdp.u2.q_esr_3_LC_2_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_3_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_3_LC_2_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_3_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13548),
            .lcout(\Lab_UT.scdp.byteToEncrypt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21100),
            .ce(N__13905),
            .sr(N__20811));
    defparam \Lab_UT.scdp.u2.q_esr_4_LC_2_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_4_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_4_LC_2_11_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_4_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__15128),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scdp.byteToEncrypt_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21100),
            .ce(N__13905),
            .sr(N__20811));
    defparam \Lab_UT.scdp.u2.q_esr_5_LC_2_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_5_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_5_LC_2_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_5_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18813),
            .lcout(\Lab_UT.scdp.byteToEncrypt_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21100),
            .ce(N__13905),
            .sr(N__20811));
    defparam \Lab_UT.scdp.u2.q_esr_6_LC_2_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_6_LC_2_11_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_6_LC_2_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_6_LC_2_11_6  (
            .in0(N__14940),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scdp.byteToEncrypt_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21100),
            .ce(N__13905),
            .sr(N__20811));
    defparam \Lab_UT.scdp.u2.q_esr_7_LC_2_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_7_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u2.q_esr_7_LC_2_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_7_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14528),
            .lcout(\Lab_UT.scdp.byteToEncrypt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21100),
            .ce(N__13905),
            .sr(N__20811));
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_3_LC_2_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_3_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_3_LC_2_12_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_3_LC_2_12_0  (
            .in0(N__9799),
            .in1(N__9854),
            .in2(N__9810),
            .in3(N__9780),
            .lcout(\Lab_UT.scdp.b2a0.N_227_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_1_7_LC_2_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_1_7_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_1_7_LC_2_12_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_1_7_LC_2_12_2  (
            .in0(N__16928),
            .in1(N__9852),
            .in2(N__9800),
            .in3(N__9778),
            .lcout(\Lab_UT.scdp.lfsrInst.N_234_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_7_LC_2_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_7_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_7_LC_2_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_7_LC_2_12_3  (
            .in0(N__9777),
            .in1(N__9792),
            .in2(N__9855),
            .in3(N__16927),
            .lcout(\Lab_UT.scdp.N_234_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_7_LC_2_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_7_LC_2_12_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_7_LC_2_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_7_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11436),
            .lcout(\Lab_UT.scdp.prng_lfsr_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21095),
            .ce(N__12792),
            .sr(N__20834));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_15_LC_2_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_15_LC_2_12_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_15_LC_2_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_15_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14154),
            .lcout(\Lab_UT.scdp.prng_lfsr_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21095),
            .ce(N__12792),
            .sr(N__20834));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_0_7_LC_2_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_0_7_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_0_7_LC_2_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNITJGS_0_7_LC_2_12_6  (
            .in0(N__16929),
            .in1(N__9853),
            .in2(N__9801),
            .in3(N__9779),
            .lcout(),
            .ltout(\Lab_UT.scdp.lfsrInst.N_234_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNILRI45_7_LC_2_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNILRI45_7_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNILRI45_7_LC_2_12_7 .LUT_INIT=16'b0011111101111111;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNILRI45_7_LC_2_12_7  (
            .in0(N__11460),
            .in1(N__11583),
            .in2(N__9765),
            .in3(N__11553),
            .lcout(\Lab_UT.scdp.g0_0_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_0_LC_2_13_0 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_2_13_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_2_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9867),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21090),
            .ce(),
            .sr(N__20837));
    defparam \buart.Z_rx.hh_1_LC_2_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_2_13_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_2_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17762),
            .lcout(buart__rx_hh_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21090),
            .ce(),
            .sr(N__20837));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_23_LC_2_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_23_LC_2_14_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_23_LC_2_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_23_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18459),
            .lcout(\Lab_UT.scdp.prng_lfsr_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21084),
            .ce(N__12791),
            .sr(N__20841));
    defparam \resetGen.shifter_ret_RNIC2S44_LC_4_3_0 .C_ON=1'b0;
    defparam \resetGen.shifter_ret_RNIC2S44_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \resetGen.shifter_ret_RNIC2S44_LC_4_3_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \resetGen.shifter_ret_RNIC2S44_LC_4_3_0  (
            .in0(N__10267),
            .in1(N__15125),
            .in2(_gnd_net_),
            .in3(N__14381),
            .lcout(\resetGen.N_421 ),
            .ltout(\resetGen.N_421_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_4_3_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_4_3_1 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \resetGen.reset_count_0_LC_4_3_1  (
            .in0(N__22561),
            .in1(_gnd_net_),
            .in2(N__9834),
            .in3(N__10181),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21142),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_4_0_o2_2_4_LC_4_3_2 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_0_o2_2_4_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.shifter_4_0_o2_2_4_LC_4_3_2 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \buart.Z_tx.shifter_4_0_o2_2_4_LC_4_3_2  (
            .in0(N__10268),
            .in1(N__15126),
            .in2(N__10206),
            .in3(N__14382),
            .lcout(\buart.Z_tx.N_554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_4_3_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_4_3_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_4_3_3 .LUT_INIT=16'b0000000010110100;
    LogicCell40 \resetGen.reset_count_1_LC_4_3_3  (
            .in0(N__22562),
            .in1(N__10182),
            .in2(N__10167),
            .in3(N__10444),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21142),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNO_0_2_LC_4_3_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_2_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_2_LC_4_3_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \resetGen.reset_count_RNO_0_2_LC_4_3_4  (
            .in0(N__10180),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10163),
            .lcout(),
            .ltout(\resetGen.N_267_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_4_3_5 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_4_3_5 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_4_3_5 .LUT_INIT=16'b0000000011001001;
    LogicCell40 \resetGen.reset_count_2_LC_4_3_5  (
            .in0(N__22563),
            .in1(N__10152),
            .in2(N__9813),
            .in3(N__10445),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21142),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNITEEC1_2_LC_4_3_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNITEEC1_2_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNITEEC1_2_LC_4_3_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \resetGen.reset_count_RNITEEC1_2_LC_4_3_6  (
            .in0(N__10179),
            .in1(N__10162),
            .in2(_gnd_net_),
            .in3(N__10151),
            .lcout(\resetGen.N_274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.tx_fsm.cstate_3_LC_4_3_7 .C_ON=1'b0;
    defparam \ufifo.tx_fsm.cstate_3_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \ufifo.tx_fsm.cstate_3_LC_4_3_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ufifo.tx_fsm.cstate_3_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(N__10135),
            .in2(_gnd_net_),
            .in3(N__15458),
            .lcout(ufifo_fifo_txdata_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21142),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.rdaddr_0_LC_4_4_0 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_0_LC_4_4_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_0_LC_4_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_0_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__10075),
            .in2(N__10139),
            .in3(N__10134),
            .lcout(\ufifo.fifo.rdaddrZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_4_0_),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_0 ),
            .clk(N__21136),
            .ce(),
            .sr(N__20818));
    defparam \ufifo.fifo.rdaddr_1_LC_4_4_1 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_1_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_1_LC_4_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_1_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(N__10042),
            .in2(_gnd_net_),
            .in3(N__10026),
            .lcout(\ufifo.fifo.rdaddrZ0Z_1 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_0 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_1 ),
            .clk(N__21136),
            .ce(),
            .sr(N__20818));
    defparam \ufifo.fifo.rdaddr_2_LC_4_4_2 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_2_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_2_LC_4_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_2_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(N__10012),
            .in2(_gnd_net_),
            .in3(N__9993),
            .lcout(\ufifo.fifo.rdaddrZ0Z_2 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_1 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_2 ),
            .clk(N__21136),
            .ce(),
            .sr(N__20818));
    defparam \ufifo.fifo.rdaddr_3_LC_4_4_3 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_3_LC_4_4_3 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_3_LC_4_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_3_LC_4_4_3  (
            .in0(_gnd_net_),
            .in1(N__9979),
            .in2(_gnd_net_),
            .in3(N__9960),
            .lcout(\ufifo.fifo.rdaddrZ0Z_3 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_2 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_3 ),
            .clk(N__21136),
            .ce(),
            .sr(N__20818));
    defparam \ufifo.fifo.rdaddr_4_LC_4_4_4 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_4_LC_4_4_4 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_4_LC_4_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_4_LC_4_4_4  (
            .in0(_gnd_net_),
            .in1(N__9946),
            .in2(_gnd_net_),
            .in3(N__9930),
            .lcout(\ufifo.fifo.rdaddrZ0Z_4 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_3 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_4 ),
            .clk(N__21136),
            .ce(),
            .sr(N__20818));
    defparam \ufifo.fifo.rdaddr_5_LC_4_4_5 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_5_LC_4_4_5 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_5_LC_4_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_5_LC_4_4_5  (
            .in0(_gnd_net_),
            .in1(N__9919),
            .in2(_gnd_net_),
            .in3(N__9900),
            .lcout(\ufifo.fifo.rdaddrZ0Z_5 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_4 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_5 ),
            .clk(N__21136),
            .ce(),
            .sr(N__20818));
    defparam \ufifo.fifo.rdaddr_6_LC_4_4_6 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_6_LC_4_4_6 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_6_LC_4_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_6_LC_4_4_6  (
            .in0(_gnd_net_),
            .in1(N__9886),
            .in2(_gnd_net_),
            .in3(N__10329),
            .lcout(\ufifo.fifo.rdaddrZ0Z_6 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_5 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_6 ),
            .clk(N__21136),
            .ce(),
            .sr(N__20818));
    defparam \ufifo.fifo.rdaddr_7_LC_4_4_7 .C_ON=1'b1;
    defparam \ufifo.fifo.rdaddr_7_LC_4_4_7 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_7_LC_4_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ufifo.fifo.rdaddr_7_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(N__10321),
            .in2(_gnd_net_),
            .in3(N__10299),
            .lcout(\ufifo.fifo.rdaddrZ0Z_7 ),
            .ltout(),
            .carryin(\ufifo.fifo.un1_rdaddr_cry_6 ),
            .carryout(\ufifo.fifo.un1_rdaddr_cry_7 ),
            .clk(N__21136),
            .ce(),
            .sr(N__20818));
    defparam \ufifo.fifo.rdaddr_8_LC_4_5_0 .C_ON=1'b0;
    defparam \ufifo.fifo.rdaddr_8_LC_4_5_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.fifo.rdaddr_8_LC_4_5_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ufifo.fifo.rdaddr_8_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(N__10288),
            .in2(_gnd_net_),
            .in3(N__10296),
            .lcout(\ufifo.fifo.rdaddrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21127),
            .ce(),
            .sr(N__20815));
    defparam \resetGen.shifter_ret_RNITHBO1_LC_4_6_0 .C_ON=1'b0;
    defparam \resetGen.shifter_ret_RNITHBO1_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \resetGen.shifter_ret_RNITHBO1_LC_4_6_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \resetGen.shifter_ret_RNITHBO1_LC_4_6_0  (
            .in0(N__13010),
            .in1(N__11130),
            .in2(N__17190),
            .in3(N__17022),
            .lcout(N_251),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_esr_2_LC_4_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_esr_2_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u0.q_esr_2_LC_4_6_1 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \Lab_UT.scdp.u0.q_esr_2_LC_4_6_1  (
            .in0(N__17023),
            .in1(N__17160),
            .in2(N__13038),
            .in3(N__16642),
            .lcout(\Lab_UT.scdp.u0.byteToDecrypt_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21122),
            .ce(N__16410),
            .sr(N__20814));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIKRN11_LC_4_6_3 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIKRN11_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIKRN11_LC_4_6_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNIKRN11_LC_4_6_3  (
            .in0(N__10245),
            .in1(N__10405),
            .in2(_gnd_net_),
            .in3(N__17159),
            .lcout(\ufifo.sb_ram512x8_inst_RNIKRN11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_4_0_o2_3_4_LC_4_6_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_0_o2_3_4_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.shifter_4_0_o2_3_4_LC_4_6_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \buart.Z_tx.shifter_4_0_o2_3_4_LC_4_6_6  (
            .in0(N__10404),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10223),
            .lcout(\buart.Z_tx.N_278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_4_7_0 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_4_7_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_4_7_0 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \resetGen.reset_count_4_LC_4_7_0  (
            .in0(N__22539),
            .in1(N__10464),
            .in2(N__10431),
            .in3(N__10452),
            .lcout(rst_ii),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21117),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.state_1_ret_LC_4_7_1 .C_ON=1'b0;
    defparam \resetGen.state_1_ret_LC_4_7_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.state_1_ret_LC_4_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \resetGen.state_1_ret_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22541),
            .lcout(rst_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21117),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_4_7_2 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_4_7_2 .LUT_INIT=16'b0000000011100001;
    LogicCell40 \resetGen.reset_count_3_LC_4_7_2  (
            .in0(N__22538),
            .in1(N__10463),
            .in2(N__10430),
            .in3(N__10451),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21117),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIKTQ21_LC_4_7_3 .C_ON=1'b0;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIKTQ21_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \ufifo.fifo.sb_ram512x8_inst_RNIKTQ21_LC_4_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ufifo.fifo.sb_ram512x8_inst_RNIKTQ21_LC_4_7_3  (
            .in0(N__10416),
            .in1(N__10356),
            .in2(_gnd_net_),
            .in3(N__16562),
            .lcout(\ufifo.sb_ram512x8_inst_RNIKTQ21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_1_iso_LC_4_7_5 .C_ON=1'b0;
    defparam \resetGen.rst_1_iso_LC_4_7_5 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_1_iso_LC_4_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_1_iso_LC_4_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22540),
            .lcout(resetGen_rst_1_iso),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21117),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_3_LC_4_7_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_3_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_3_LC_4_7_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_3_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(N__17735),
            .in2(_gnd_net_),
            .in3(N__14909),
            .lcout(N_233_reti),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI679E_6_LC_4_7_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI679E_6_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI679E_6_LC_4_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNI679E_6_LC_4_7_7  (
            .in0(N__10665),
            .in1(N__10491),
            .in2(_gnd_net_),
            .in3(N__10836),
            .lcout(\Lab_UT.scdp.msBitsi.q_esr_RNI679EZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lsBitsi.q_esr_2_LC_4_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_2_LC_4_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_2_LC_4_8_0 .LUT_INIT=16'b0000111011100000;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_esr_2_LC_4_8_0  (
            .in0(N__10539),
            .in1(N__10556),
            .in2(N__10590),
            .in3(N__12638),
            .lcout(\Lab_UT.scdp.lsBitsD_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21110),
            .ce(N__11217),
            .sr(N__20809));
    defparam \Lab_UT.scdp.lsBitsi.q_esr_4_LC_4_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_4_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_4_LC_4_8_1 .LUT_INIT=16'b0000100111111111;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_esr_4_LC_4_8_1  (
            .in0(N__12639),
            .in1(N__10588),
            .in2(N__10560),
            .in3(N__11693),
            .lcout(\Lab_UT.scdp.lsBitsD_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21110),
            .ce(N__11217),
            .sr(N__20809));
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_o2_2_LC_4_8_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_o2_2_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_o2_2_LC_4_8_2 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \Lab_UT.scdp.b2a1.asciiHex_2_i_o2_2_LC_4_8_2  (
            .in0(N__11691),
            .in1(N__10343),
            .in2(_gnd_net_),
            .in3(N__12707),
            .lcout(\Lab_UT.scdp.b2a1.N_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lsBitsi.q_esr_0_LC_4_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_0_LC_4_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_0_LC_4_8_3 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_esr_0_LC_4_8_3  (
            .in0(N__12708),
            .in1(N__10476),
            .in2(N__10347),
            .in3(N__11692),
            .lcout(\Lab_UT.scdp.lsBitsD_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21110),
            .ce(N__11217),
            .sr(N__20809));
    defparam \Lab_UT.scdp.b2a1.lsBits_i_0_o2_6_LC_4_8_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a1.lsBits_i_0_o2_6_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a1.lsBits_i_0_o2_6_LC_4_8_4 .LUT_INIT=16'b0111010101010111;
    LogicCell40 \Lab_UT.scdp.b2a1.lsBits_i_0_o2_6_LC_4_8_4  (
            .in0(N__11690),
            .in1(N__10554),
            .in2(N__10589),
            .in3(N__12636),
            .lcout(\Lab_UT.scdp.lsBits_i_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_x2_0_2_LC_4_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_x2_0_2_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_x2_0_2_LC_4_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.scdp.b2a1.asciiHex_2_i_x2_0_2_LC_4_8_5  (
            .in0(N__10602),
            .in1(N__11847),
            .in2(_gnd_net_),
            .in3(N__11660),
            .lcout(\Lab_UT.scdp.b2a1.N_220_i ),
            .ltout(\Lab_UT.scdp.b2a1.N_220_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_o2_3_LC_4_8_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_o2_3_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_o2_3_LC_4_8_6 .LUT_INIT=16'b1111010111111010;
    LogicCell40 \Lab_UT.scdp.b2a1.asciiHex_2_i_o2_3_LC_4_8_6  (
            .in0(N__10584),
            .in1(_gnd_net_),
            .in2(N__10563),
            .in3(N__12637),
            .lcout(\Lab_UT.scdp.N_282 ),
            .ltout(\Lab_UT.scdp.N_282_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lsBitsi.q_esr_1_LC_4_8_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_1_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_esr_1_LC_4_8_7 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_esr_1_LC_4_8_7  (
            .in0(N__10555),
            .in1(_gnd_net_),
            .in2(N__10542),
            .in3(N__10538),
            .lcout(\Lab_UT.scdp.lsBitsD_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21110),
            .ce(N__11217),
            .sr(N__20809));
    defparam \Lab_UT.scctrl.state_1_ret_5_RNI1UBG9_LC_4_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNI1UBG9_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNI1UBG9_LC_4_9_1 .LUT_INIT=16'b0000010000001110;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_5_RNI1UBG9_LC_4_9_1  (
            .in0(N__11346),
            .in1(N__10526),
            .in2(N__20141),
            .in3(N__14000),
            .lcout(\Lab_UT.scctrl.sccLdLFSR ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lsBitsi.q_5_LC_4_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_5_LC_4_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_5_LC_4_9_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_5_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(N__10862),
            .in2(_gnd_net_),
            .in3(N__11231),
            .lcout(\Lab_UT.scdp.lsBitsi.lsBitsDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21101),
            .ce(),
            .sr(N__20812));
    defparam \Lab_UT.scctrl.state_ret_13_RNI7RC32_LC_4_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNI7RC32_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNI7RC32_LC_4_9_3 .LUT_INIT=16'b0100010101000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNI7RC32_LC_4_9_3  (
            .in0(N__20114),
            .in1(N__10509),
            .in2(N__21723),
            .in3(N__23127),
            .lcout(\Lab_UT.scctrl.EmsLoaded ),
            .ltout(\Lab_UT.scctrl.EmsLoaded_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNICOE1_0_LC_4_9_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNICOE1_0_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNICOE1_0_LC_4_9_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNICOE1_0_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10503),
            .in3(N__21706),
            .lcout(\Lab_UT.sccElsBitsLd ),
            .ltout(\Lab_UT.sccElsBitsLd_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lsBitsi.q_6_LC_4_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_6_LC_4_9_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_6_LC_4_9_5 .LUT_INIT=16'b0000110011111100;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_6_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(N__10490),
            .in2(N__10500),
            .in3(N__10497),
            .lcout(\Lab_UT.scdp.lsBitsD_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21101),
            .ce(),
            .sr(N__20812));
    defparam \Lab_UT.scdp.lsBitsi.q_3_LC_4_9_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lsBitsi.q_3_LC_4_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.lsBitsi.q_3_LC_4_9_7 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \Lab_UT.scdp.lsBitsi.q_3_LC_4_9_7  (
            .in0(N__11232),
            .in1(N__10787),
            .in2(N__11697),
            .in3(N__10475),
            .lcout(\Lab_UT.scdp.lsBitsD_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21101),
            .ce(),
            .sr(N__20812));
    defparam \Lab_UT.scdp.msBitsi.q_esr_1_LC_4_10_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_1_LC_4_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_1_LC_4_10_0 .LUT_INIT=16'b1010101010011000;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_1_LC_4_10_0  (
            .in0(N__10630),
            .in1(N__10693),
            .in2(N__10724),
            .in3(N__11870),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsD_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21096),
            .ce(N__11216),
            .sr(N__20813));
    defparam \Lab_UT.scdp.msBitsi.q_esr_0_LC_4_10_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_0_LC_4_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_0_LC_4_10_1 .LUT_INIT=16'b1010010110100110;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_0_LC_4_10_1  (
            .in0(N__11869),
            .in1(N__10715),
            .in2(N__10700),
            .in3(N__10629),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsD_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21096),
            .ce(N__11216),
            .sr(N__20813));
    defparam \Lab_UT.scdp.msBitsi.q_esr_2_LC_4_10_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_2_LC_4_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_2_LC_4_10_2 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_2_LC_4_10_2  (
            .in0(N__10631),
            .in1(N__10694),
            .in2(N__10725),
            .in3(N__11871),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsD_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21096),
            .ce(N__11216),
            .sr(N__20813));
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_1_1_LC_4_10_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_1_1_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_1_1_LC_4_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_1_1_LC_4_10_3  (
            .in0(N__11059),
            .in1(N__12570),
            .in2(N__10743),
            .in3(N__11079),
            .lcout(\Lab_UT.scdp.b2a0.N_238_i ),
            .ltout(\Lab_UT.scdp.b2a0.N_238_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_4_LC_4_10_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_4_LC_4_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_4_LC_4_10_4 .LUT_INIT=16'b1010111010101011;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_4_LC_4_10_4  (
            .in0(N__10696),
            .in1(N__10653),
            .in2(N__10728),
            .in3(N__11976),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsD_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21096),
            .ce(N__11216),
            .sr(N__20813));
    defparam \Lab_UT.scdp.msBitsi.q_esr_3_LC_4_10_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_3_LC_4_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_3_LC_4_10_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_3_LC_4_10_5  (
            .in0(N__10695),
            .in1(N__10722),
            .in2(_gnd_net_),
            .in3(N__10632),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsD_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21096),
            .ce(N__11216),
            .sr(N__20813));
    defparam \Lab_UT.scdp.msBitsi.q_esr_6_LC_4_10_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_6_LC_4_10_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_6_LC_4_10_6 .LUT_INIT=16'b0000101100001110;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_6_LC_4_10_6  (
            .in0(N__10723),
            .in1(N__10652),
            .in2(N__10701),
            .in3(N__11975),
            .lcout(\Lab_UT.scdp.msBitsi.msBitsD_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21096),
            .ce(N__11216),
            .sr(N__20813));
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_0_1_LC_4_10_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_0_1_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_0_1_LC_4_10_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.scdp.b2a0.asciiHex_2_i_x2_0_1_LC_4_10_7  (
            .in0(N__11974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10651),
            .lcout(\Lab_UT.scdp.b2a0.N_224_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI3LL8_0_LC_4_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI3LL8_0_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI3LL8_0_LC_4_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNI3LL8_0_LC_4_11_0  (
            .in0(N__10617),
            .in1(N__10611),
            .in2(_gnd_net_),
            .in3(N__10828),
            .lcout(\Lab_UT.scdp.msBitsi.N_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8_1_LC_4_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8_1_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8_1_LC_4_11_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNI5NL8_1_LC_4_11_1  (
            .in0(N__10829),
            .in1(N__10932),
            .in2(_gnd_net_),
            .in3(N__10926),
            .lcout(),
            .ltout(\Lab_UT.scdp.msBitsi.N_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_1_LC_4_11_2 .C_ON=1'b0;
    defparam \ufifo.txdataD_1_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_1_LC_4_11_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ufifo.txdataD_1_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__21709),
            .in2(N__10917),
            .in3(N__10974),
            .lcout(\ufifo.txdataDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21091),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI7PL8_2_LC_4_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI7PL8_2_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI7PL8_2_LC_4_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNI7PL8_2_LC_4_11_3  (
            .in0(N__10831),
            .in1(N__10902),
            .in2(_gnd_net_),
            .in3(N__10896),
            .lcout(\Lab_UT.scdp.msBitsi.N_1919_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNIBTL8_4_LC_4_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNIBTL8_4_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNIBTL8_4_LC_4_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNIBTL8_4_LC_4_11_4  (
            .in0(N__10884),
            .in1(N__10878),
            .in2(_gnd_net_),
            .in3(N__10832),
            .lcout(\Lab_UT.scdp.msBitsi.N_1917_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNI2JO42_1_LC_4_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNI2JO42_1_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNI2JO42_1_LC_4_11_5 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \Lab_UT.scdp.u0.q_RNI2JO42_1_LC_4_11_5  (
            .in0(N__12088),
            .in1(N__12034),
            .in2(_gnd_net_),
            .in3(N__11971),
            .lcout(),
            .ltout(\Lab_UT.scdp.N_332_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_5_LC_4_11_6 .C_ON=1'b0;
    defparam \ufifo.txdataD_5_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_5_LC_4_11_6 .LUT_INIT=16'b1110001011101110;
    LogicCell40 \ufifo.txdataD_5_LC_4_11_6  (
            .in0(N__10869),
            .in1(N__21710),
            .in2(N__10851),
            .in3(N__11552),
            .lcout(\ufifo.txdataDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21091),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI019E_3_LC_4_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI019E_3_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_RNI019E_3_LC_4_11_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_RNI019E_3_LC_4_11_7  (
            .in0(N__10830),
            .in1(_gnd_net_),
            .in2(N__10797),
            .in3(N__10788),
            .lcout(\Lab_UT.scdp.msBitsi.N_1915_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_3_LC_4_12_0 .C_ON=1'b0;
    defparam \ufifo.txdataD_3_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_3_LC_4_12_0 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \ufifo.txdataD_3_LC_4_12_0  (
            .in0(N__10773),
            .in1(N__10764),
            .in2(N__21729),
            .in3(N__11085),
            .lcout(\ufifo.txdataDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21085),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_2_LC_4_12_1 .C_ON=1'b0;
    defparam \ufifo.txdataD_2_LC_4_12_1 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_2_LC_4_12_1 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \ufifo.txdataD_2_LC_4_12_1  (
            .in0(N__21707),
            .in1(N__11922),
            .in2(N__11022),
            .in3(N__11736),
            .lcout(\ufifo.txdataDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21085),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_4_LC_4_12_2 .C_ON=1'b0;
    defparam \ufifo.txdataD_4_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_4_LC_4_12_2 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \ufifo.txdataD_4_LC_4_12_2  (
            .in0(N__10941),
            .in1(N__21708),
            .in2(N__10998),
            .in3(N__11094),
            .lcout(\ufifo.txdataDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21085),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNI4GMQ4_1_LC_4_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNI4GMQ4_1_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNI4GMQ4_1_LC_4_12_3 .LUT_INIT=16'b1111111110010110;
    LogicCell40 \Lab_UT.scdp.u1.q_RNI4GMQ4_1_LC_4_12_3  (
            .in0(N__11846),
            .in1(N__11656),
            .in2(N__11628),
            .in3(N__11384),
            .lcout(\Lab_UT.scdp.N_552 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_esr_RNIA29D1_0_2_LC_4_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_esr_RNIA29D1_0_2_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_esr_RNIA29D1_0_2_LC_4_12_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.u0.q_esr_RNIA29D1_0_2_LC_4_12_4  (
            .in0(N__12568),
            .in1(N__10965),
            .in2(N__11060),
            .in3(N__11074),
            .lcout(\Lab_UT.scdp.N_228_i_0 ),
            .ltout(\Lab_UT.scdp.N_228_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNI2TTL2_1_LC_4_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNI2TTL2_1_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNI2TTL2_1_LC_4_12_5 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNI2TTL2_1_LC_4_12_5  (
            .in0(N__11623),
            .in1(N__11845),
            .in2(N__10968),
            .in3(N__11655),
            .lcout(\Lab_UT.scdp.u1.g0_0_i_a5_0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_esr_RNIA29D1_2_LC_4_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_esr_RNIA29D1_2_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_esr_RNIA29D1_2_LC_4_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.u0.q_esr_RNIA29D1_2_LC_4_12_6  (
            .in0(N__12569),
            .in1(N__10964),
            .in2(N__11061),
            .in3(N__11075),
            .lcout(\Lab_UT.scdp.N_228_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNI5V781_0_1_LC_4_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNI5V781_0_1_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNI5V781_0_1_LC_4_12_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.scdp.u0.q_RNI5V781_0_1_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(N__12022),
            .in2(_gnd_net_),
            .in3(N__11955),
            .lcout(\Lab_UT.scdp.N_225_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNICF9Q4_7_LC_4_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNICF9Q4_7_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNICF9Q4_7_LC_4_13_0 .LUT_INIT=16'b0011011111111111;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNICF9Q4_7_LC_4_13_0  (
            .in0(N__11546),
            .in1(N__10953),
            .in2(N__11109),
            .in3(N__11792),
            .lcout(\Lab_UT.scdp.g0_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIPUDN_17_LC_4_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIPUDN_17_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIPUDN_17_LC_4_13_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIPUDN_17_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__11142),
            .in2(_gnd_net_),
            .in3(N__11034),
            .lcout(\Lab_UT.scdp.d2eData_3_0_1 ),
            .ltout(\Lab_UT.scdp.d2eData_3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNI116R2_1_LC_4_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNI116R2_1_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNI116R2_1_LC_4_13_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNI116R2_1_LC_4_13_2  (
            .in0(N__11575),
            .in1(N__11621),
            .in2(N__10935),
            .in3(N__11840),
            .lcout(),
            .ltout(\Lab_UT.scdp.u1.g0_0_i_a5_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNI7PSB8_0_LC_4_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNI7PSB8_0_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNI7PSB8_0_LC_4_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNI7PSB8_0_LC_4_13_3  (
            .in0(N__12717),
            .in1(N__11108),
            .in2(N__11097),
            .in3(N__11547),
            .lcout(\Lab_UT.scdp.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNIOKSG2_1_LC_4_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNIOKSG2_1_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNIOKSG2_1_LC_4_13_4 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNIOKSG2_1_LC_4_13_4  (
            .in0(N__11841),
            .in1(N__11791),
            .in2(N__11661),
            .in3(N__11622),
            .lcout(),
            .ltout(\Lab_UT.scdp.u1.g0_0_i_a5_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNIUCJ18_0_LC_4_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNIUCJ18_0_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNIUCJ18_0_LC_4_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNIUCJ18_0_LC_4_13_5  (
            .in0(N__12600),
            .in1(N__11459),
            .in2(N__11088),
            .in3(N__11548),
            .lcout(\Lab_UT.scdp.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIHOFN_22_LC_4_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIHOFN_22_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIHOFN_22_LC_4_13_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIHOFN_22_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__11136),
            .in2(_gnd_net_),
            .in3(N__11028),
            .lcout(\Lab_UT.scdp.d2eData_3_0_a2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNICL1I3_1_LC_4_13_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNICL1I3_1_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNICL1I3_1_LC_4_13_7 .LUT_INIT=16'b0011001110110111;
    LogicCell40 \Lab_UT.scdp.u0.q_RNICL1I3_1_LC_4_13_7  (
            .in0(N__11963),
            .in1(N__12089),
            .in2(N__12048),
            .in3(N__11545),
            .lcout(\Lab_UT.scdp.N_276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_1_LC_4_14_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_1_LC_4_14_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_1_LC_4_14_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_1_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__17526),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21077),
            .ce(N__12788),
            .sr(N__20850));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_14_LC_4_14_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_14_LC_4_14_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_14_LC_4_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_14_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13926),
            .lcout(\Lab_UT.scdp.prng_lfsr_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21077),
            .ce(N__12788),
            .sr(N__20850));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_17_LC_4_14_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_17_LC_4_14_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_17_LC_4_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_17_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16890),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21077),
            .ce(N__12788),
            .sr(N__20850));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_22_LC_4_14_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_22_LC_4_14_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_22_LC_4_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_22_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14103),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21077),
            .ce(N__12788),
            .sr(N__20850));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_25_LC_4_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_25_LC_4_14_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_25_LC_4_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_25_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16851),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21077),
            .ce(N__12788),
            .sr(N__20850));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_3_LC_4_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_3_LC_4_14_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_3_LC_4_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_3_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11415),
            .lcout(\Lab_UT.scdp.prng_lfsr_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21077),
            .ce(N__12788),
            .sr(N__20850));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_30_LC_4_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_30_LC_4_14_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_30_LC_4_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_30_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12501),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21077),
            .ce(N__12788),
            .sr(N__20850));
    defparam \Lab_UT.scctrl.state_1_RNO_9_0_LC_5_3_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_9_0_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_9_0_LC_5_3_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_9_0_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__13223),
            .in2(_gnd_net_),
            .in3(N__22058),
            .lcout(\Lab_UT.scctrl.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.val_0_a2_3_3_LC_5_3_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_0_a2_3_3_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_0_a2_3_3_LC_5_3_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.scdp.a2b.val_0_a2_3_3_LC_5_3_6  (
            .in0(N__13541),
            .in1(N__17162),
            .in2(_gnd_net_),
            .in3(N__13031),
            .lcout(\Lab_UT.N_540i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.shifter_ret_LC_5_4_7 .C_ON=1'b0;
    defparam \resetGen.shifter_ret_LC_5_4_7 .SEQ_MODE=4'b1011;
    defparam \resetGen.shifter_ret_LC_5_4_7 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \resetGen.shifter_ret_LC_5_4_7  (
            .in0(N__11253),
            .in1(N__14526),
            .in2(_gnd_net_),
            .in3(N__15116),
            .lcout(\resetGen.N_243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21128),
            .ce(N__13448),
            .sr(N__20848));
    defparam \buart.Z_rx.shifter_ret_2_LC_5_5_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_2_LC_5_5_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_2_LC_5_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_2_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18780),
            .lcout(\buart.bu_rx_data_i_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21123),
            .ce(N__13446),
            .sr(N__20842));
    defparam \Lab_UT.scctrl.shifter_ret_6_LC_5_5_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_6_LC_5_5_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.shifter_ret_6_LC_5_5_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_6_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(N__18781),
            .in2(_gnd_net_),
            .in3(N__15084),
            .lcout(\Lab_UT.scctrl.N_534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21123),
            .ce(N__13446),
            .sr(N__20842));
    defparam \buart.Z_rx.shifter_1_5_LC_5_5_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_5_LC_5_5_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_5_LC_5_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_5_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14900),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21123),
            .ce(N__13446),
            .sr(N__20842));
    defparam \buart.Z_rx.shifter_2_6_LC_5_5_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_6_LC_5_5_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_6_LC_5_5_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_2_6_LC_5_5_7  (
            .in0(N__14527),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21123),
            .ce(N__13446),
            .sr(N__20842));
    defparam \Lab_UT.scctrl.next_state_1_i_i_o2_5_0_LC_5_6_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_1_i_i_o2_5_0_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_1_i_i_o2_5_0_LC_5_6_0 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \Lab_UT.scctrl.next_state_1_i_i_o2_5_0_LC_5_6_0  (
            .in0(N__13501),
            .in1(N__17161),
            .in2(_gnd_net_),
            .in3(N__15075),
            .lcout(\Lab_UT.scctrl.N_259i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_6_LC_5_6_1 .C_ON=1'b0;
    defparam \ufifo.txdataD_6_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_6_LC_5_6_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ufifo.txdataD_6_LC_5_6_1  (
            .in0(N__11193),
            .in1(N__21721),
            .in2(_gnd_net_),
            .in3(N__11514),
            .lcout(\ufifo.txdataDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21118),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_5_RNIOMGF_LC_5_6_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_5_RNIOMGF_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_5_RNIOMGF_LC_5_6_4 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_5_RNIOMGF_LC_5_6_4  (
            .in0(N__18755),
            .in1(N__11172),
            .in2(_gnd_net_),
            .in3(N__12171),
            .lcout(\Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0 ),
            .ltout(\Lab_UT.scctrl.next_state_1_i_i_o2_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_1_RNI4BLT2_LC_5_6_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_1_RNI4BLT2_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_1_RNI4BLT2_LC_5_6_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scctrl.state_ret_1_RNI4BLT2_LC_5_6_5  (
            .in0(N__18275),
            .in1(N__14522),
            .in2(N__11166),
            .in3(N__14380),
            .lcout(\Lab_UT.scctrl.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_9_LC_5_6_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_9_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_9_LC_5_6_6 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_9_LC_5_6_6  (
            .in0(N__22043),
            .in1(N__19731),
            .in2(N__22441),
            .in3(N__22292),
            .lcout(\Lab_UT.scctrl.N_415_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_8_LC_5_6_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_8_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_8_LC_5_6_7 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_8_LC_5_6_7  (
            .in0(N__22820),
            .in1(N__18065),
            .in2(N__15430),
            .in3(N__14632),
            .lcout(\Lab_UT.scctrl.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_4_LC_5_7_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_4_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_4_LC_5_7_1 .LUT_INIT=16'b0100000001010000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_4_LC_5_7_1  (
            .in0(N__11163),
            .in1(N__23202),
            .in2(N__11157),
            .in3(N__22970),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g1_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_1_LC_5_7_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_1_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_1_LC_5_7_2 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_1_LC_5_7_2  (
            .in0(N__12129),
            .in1(N__23690),
            .in2(N__11148),
            .in3(N__23507),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_LC_5_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_ret_2_LC_5_7_3 .LUT_INIT=16'b0000001010101010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_LC_5_7_3  (
            .in0(N__22542),
            .in1(N__14742),
            .in2(N__11145),
            .in3(N__15398),
            .lcout(\Lab_UT.scctrl.N_351_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21111),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txDataValidD_LC_5_7_4 .C_ON=1'b0;
    defparam \ufifo.txDataValidD_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \ufifo.txDataValidD_LC_5_7_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ufifo.txDataValidD_LC_5_7_4  (
            .in0(N__13614),
            .in1(N__11493),
            .in2(_gnd_net_),
            .in3(N__13626),
            .lcout(\ufifo.txDataValidDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21111),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.un3_reset_count_i_o2_3_LC_5_7_7 .C_ON=1'b0;
    defparam \resetGen.un3_reset_count_i_o2_3_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \resetGen.un3_reset_count_i_o2_3_LC_5_7_7 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \resetGen.un3_reset_count_i_o2_3_LC_5_7_7  (
            .in0(N__11249),
            .in1(N__14468),
            .in2(_gnd_net_),
            .in3(N__15079),
            .lcout(N_243_reti),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_0_RNIQM5P_LC_5_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_0_RNIQM5P_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_0_RNIQM5P_LC_5_8_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_0_RNIQM5P_LC_5_8_0  (
            .in0(N__12974),
            .in1(N__13144),
            .in2(_gnd_net_),
            .in3(N__13170),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g1_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_0_RNIK3S32_LC_5_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_0_RNIK3S32_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_0_RNIK3S32_LC_5_8_1 .LUT_INIT=16'b1010101001000000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_0_RNIK3S32_LC_5_8_1  (
            .in0(N__15104),
            .in1(N__17827),
            .in2(N__11235),
            .in3(N__15180),
            .lcout(\Lab_UT.scctrl.g1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_fast_1_LC_5_8_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_1_LC_5_8_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_1_LC_5_8_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_fast_1_LC_5_8_4  (
            .in0(N__12975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buart__rx_shifter_0_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21102),
            .ce(N__13441),
            .sr(N__20830));
    defparam \buart.Z_rx.shifter_0_1_LC_5_8_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_1_LC_5_8_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_1_LC_5_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_1_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12976),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21102),
            .ce(N__13441),
            .sr(N__20830));
    defparam \Lab_UT.scctrl.shifter_ret_0_LC_5_8_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_0_LC_5_8_6 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.scctrl.shifter_ret_0_LC_5_8_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_0_LC_5_8_6  (
            .in0(N__13508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17155),
            .lcout(\Lab_UT.scctrl.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21102),
            .ce(N__13441),
            .sr(N__20830));
    defparam \buart.Z_rx.shifter_0_2_LC_5_8_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_2_LC_5_8_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_2_LC_5_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_2_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13509),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21102),
            .ce(N__13441),
            .sr(N__20830));
    defparam \Lab_UT.scdp.msBitsi.q_esr_ctle_6_LC_5_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.msBitsi.q_esr_ctle_6_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.msBitsi.q_esr_ctle_6_LC_5_9_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scdp.msBitsi.q_esr_ctle_6_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__16447),
            .in2(_gnd_net_),
            .in3(N__11230),
            .lcout(\Lab_UT.scdp.sccElsBitsLd_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_0_RNIDPMQ_LC_5_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_0_RNIDPMQ_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_0_RNIDPMQ_LC_5_9_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_0_RNIDPMQ_LC_5_9_2  (
            .in0(N__17128),
            .in1(N__12983),
            .in2(_gnd_net_),
            .in3(N__13171),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_0_RNI76D52_LC_5_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_0_RNI76D52_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_0_RNI76D52_LC_5_9_3 .LUT_INIT=16'b1100110000100000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_0_RNI76D52_LC_5_9_3  (
            .in0(N__17855),
            .in1(N__15183),
            .in2(N__11394),
            .in3(N__15124),
            .lcout(\Lab_UT.scctrl.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_1_LC_5_9_4 .C_ON=1'b0;
    defparam \resetGen.rst_1_LC_5_9_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_1_LC_5_9_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \resetGen.rst_1_LC_5_9_4  (
            .in0(N__22548),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21097),
            .ce(),
            .sr(_gnd_net_));
    defparam \ufifo.txdataD_0_LC_5_9_5 .C_ON=1'b0;
    defparam \ufifo.txdataD_0_LC_5_9_5 .SEQ_MODE=4'b1000;
    defparam \ufifo.txdataD_0_LC_5_9_5 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \ufifo.txdataD_0_LC_5_9_5  (
            .in0(N__21724),
            .in1(N__11391),
            .in2(N__11373),
            .in3(N__12735),
            .lcout(\ufifo.txdataDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21097),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_5_RNIDAO06_LC_5_9_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNIDAO06_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNIDAO06_LC_5_9_6 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_5_RNIDAO06_LC_5_9_6  (
            .in0(N__23126),
            .in1(N__18278),
            .in2(N__20328),
            .in3(N__13984),
            .lcout(\Lab_UT.scctrl.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIJOOS_LC_5_9_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIJOOS_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIJOOS_LC_5_9_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNIJOOS_LC_5_9_7  (
            .in0(N__20664),
            .in1(N__20118),
            .in2(_gnd_net_),
            .in3(N__21408),
            .lcout(\Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0dup_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_4_LC_5_10_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_4_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_4_LC_5_10_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIPVCP_4_LC_5_10_0  (
            .in0(N__13668),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13724),
            .lcout(\buart.Z_rx.sample_i_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.rddataDV.q_0_LC_5_10_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.rddataDV.q_0_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.rddataDV.q_0_LC_5_10_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.scdp.rddataDV.q_0_LC_5_10_1  (
            .in0(N__13725),
            .in1(N__13669),
            .in2(N__11325),
            .in3(N__13860),
            .lcout(\Lab_UT.scdp.binVal_ValidD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21092),
            .ce(),
            .sr(N__20816));
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_2_LC_5_10_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_2_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_2_LC_5_10_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIPVCP_2_LC_5_10_2  (
            .in0(N__13792),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13821),
            .lcout(\buart.Z_rx.N_230 ),
            .ltout(\buart.Z_rx.N_230_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_5_10_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_5_10_3 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_5_10_3  (
            .in0(N__13723),
            .in1(N__13667),
            .in2(N__11439),
            .in3(N__13859),
            .lcout(N_232),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.k0h.q_2_LC_5_10_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0h.q_2_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0h.q_2_LC_5_10_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k0h.q_2_LC_5_10_4  (
            .in0(N__18574),
            .in1(N__16799),
            .in2(N__12587),
            .in3(N__12478),
            .lcout(\Lab_UT.scdp.key0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21092),
            .ce(),
            .sr(N__20816));
    defparam \Lab_UT.scdp.k0h.q_3_LC_5_10_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0h.q_3_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0h.q_3_LC_5_10_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.scdp.k0h.q_3_LC_5_10_5  (
            .in0(N__12479),
            .in1(N__18576),
            .in2(N__11432),
            .in3(N__18533),
            .lcout(\Lab_UT.scdp.key0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21092),
            .ce(),
            .sr(N__20816));
    defparam \Lab_UT.scdp.k0l.q_2_LC_5_10_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0l.q_2_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0l.q_2_LC_5_10_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k0l.q_2_LC_5_10_6  (
            .in0(N__18575),
            .in1(N__16800),
            .in2(N__11762),
            .in3(N__17555),
            .lcout(\Lab_UT.scdp.key0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21092),
            .ce(),
            .sr(N__20816));
    defparam \Lab_UT.scdp.k0l.q_3_LC_5_10_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0l.q_3_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0l.q_3_LC_5_10_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.scdp.k0l.q_3_LC_5_10_7  (
            .in0(N__17556),
            .in1(N__18534),
            .in2(N__18623),
            .in3(N__11408),
            .lcout(\Lab_UT.scdp.key0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21092),
            .ce(),
            .sr(N__20816));
    defparam \Lab_UT.scdp.rxdataD.q_1_LC_5_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.rxdataD.q_1_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.rxdataD.q_1_LC_5_11_0 .LUT_INIT=16'b1100110111001001;
    LogicCell40 \Lab_UT.scdp.rxdataD.q_1_LC_5_11_0  (
            .in0(N__17051),
            .in1(N__17166),
            .in2(N__16641),
            .in3(N__13020),
            .lcout(\Lab_UT.scdp.binValD_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21086),
            .ce(),
            .sr(N__20819));
    defparam \Lab_UT.scdp.rxdataD.q_2_LC_5_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.rxdataD.q_2_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.rxdataD.q_2_LC_5_11_1 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \Lab_UT.scdp.rxdataD.q_2_LC_5_11_1  (
            .in0(N__17165),
            .in1(N__13018),
            .in2(N__16639),
            .in3(N__17052),
            .lcout(\Lab_UT.scdp.binValD_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21086),
            .ce(),
            .sr(N__20819));
    defparam \Lab_UT.scdp.a2b.val_0_2_LC_5_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_0_2_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_0_2_LC_5_11_2 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \Lab_UT.scdp.a2b.val_0_2_LC_5_11_2  (
            .in0(N__17050),
            .in1(N__17164),
            .in2(N__16640),
            .in3(N__13019),
            .lcout(),
            .ltout(\Lab_UT.scdp.binVal_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_2_LC_5_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_2_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u1.q_2_LC_5_11_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \Lab_UT.scdp.u1.q_2_LC_5_11_3  (
            .in0(N__21593),
            .in1(N__12665),
            .in2(N__11397),
            .in3(N__21624),
            .lcout(\Lab_UT.scdp.u1.byteToDecryptZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21086),
            .ce(),
            .sr(N__20819));
    defparam \Lab_UT.scdp.u1.q_1_LC_5_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_1_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u1.q_1_LC_5_11_4 .LUT_INIT=16'b0111111100100000;
    LogicCell40 \Lab_UT.scdp.u1.q_1_LC_5_11_4  (
            .in0(N__21623),
            .in1(N__11502),
            .in2(N__21594),
            .in3(N__11617),
            .lcout(\Lab_UT.scdp.u1.byteToDecrypt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21086),
            .ce(),
            .sr(N__20819));
    defparam \Lab_UT.scdp.a2b.val_i_1_LC_5_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_i_1_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_i_1_LC_5_11_5 .LUT_INIT=16'b0101010101010010;
    LogicCell40 \Lab_UT.scdp.a2b.val_i_1_LC_5_11_5  (
            .in0(N__17163),
            .in1(N__13017),
            .in2(N__16638),
            .in3(N__17049),
            .lcout(\Lab_UT.scdp.N_73 ),
            .ltout(\Lab_UT.scdp.N_73_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_1_LC_5_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_1_LC_5_11_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u0.q_1_LC_5_11_6 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \Lab_UT.scdp.u0.q_1_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__12035),
            .in2(N__11496),
            .in3(N__16956),
            .lcout(\Lab_UT.scdp.byteToDecrypt_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21086),
            .ce(),
            .sr(N__20819));
    defparam \Lab_UT.scctrl.r5.q_0_LC_5_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.r5.q_0_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.r5.q_0_LC_5_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.r5.q_0_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__21589),
            .in2(_gnd_net_),
            .in3(N__21622),
            .lcout(\Lab_UT.scctrl.delayload ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21086),
            .ce(),
            .sr(N__20819));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_29_LC_5_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_29_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_29_LC_5_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_29_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12525),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21080),
            .ce(N__12790),
            .sr(N__20847));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_5_LC_5_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_5_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_5_LC_5_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_5_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12455),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21080),
            .ce(N__12790),
            .sr(N__20847));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_13_LC_5_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_13_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_13_LC_5_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_13_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17481),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21080),
            .ce(N__12790),
            .sr(N__20847));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIRBV41_5_LC_5_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIRBV41_5_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIRBV41_5_LC_5_12_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIRBV41_5_LC_5_12_3  (
            .in0(N__11445),
            .in1(N__11484),
            .in2(N__11478),
            .in3(N__11469),
            .lcout(\Lab_UT.scdp.d2eData_3_5 ),
            .ltout(\Lab_UT.scdp.d2eData_3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNI5V781_1_LC_5_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNI5V781_1_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNI5V781_1_LC_5_12_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \Lab_UT.scdp.u0.q_RNI5V781_1_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11463),
            .in3(N__12021),
            .lcout(\Lab_UT.scdp.N_225_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_21_LC_5_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_21_LC_5_12_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_21_LC_5_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_21_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14040),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21080),
            .ce(N__12790),
            .sr(N__20847));
    defparam \Lab_UT.scdp.u1.q_RNIOKSG2_0_LC_5_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNIOKSG2_0_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNIOKSG2_0_LC_5_12_6 .LUT_INIT=16'b0001010000101000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNIOKSG2_0_LC_5_12_6  (
            .in0(N__12698),
            .in1(N__11962),
            .in2(N__12043),
            .in3(N__17267),
            .lcout(),
            .ltout(\Lab_UT.scdp.u1.g0_0_i_a5_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNI3IJ18_0_LC_5_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNI3IJ18_0_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNI3IJ18_0_LC_5_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNI3IJ18_0_LC_5_12_7  (
            .in0(N__11579),
            .in1(N__11796),
            .in2(N__11745),
            .in3(N__11742),
            .lcout(\Lab_UT.scdp.N_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIT2EN_19_LC_5_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIT2EN_19_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIT2EN_19_LC_5_13_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIT2EN_19_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__11892),
            .in2(_gnd_net_),
            .in3(N__11667),
            .lcout(\Lab_UT.scdp.d2eData_3_0_3 ),
            .ltout(\Lab_UT.scdp.d2eData_3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI96HI1_3_LC_5_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI96HI1_3_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI96HI1_3_LC_5_13_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI96HI1_3_LC_5_13_1  (
            .in0(N__12830),
            .in1(N__11726),
            .in2(N__11730),
            .in3(N__16665),
            .lcout(\Lab_UT.scdp.N_255_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_x2_3_LC_5_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_x2_3_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a1.asciiHex_2_i_x2_3_LC_5_13_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.b2a1.asciiHex_2_i_x2_3_LC_5_13_2  (
            .in0(N__11727),
            .in1(N__12831),
            .in2(N__11718),
            .in3(N__11703),
            .lcout(\Lab_UT.scdp.N_226_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_19_LC_5_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_19_LC_5_13_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_19_LC_5_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_19_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17430),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21078),
            .ce(N__12789),
            .sr(N__20851));
    defparam \Lab_UT.scdp.u1.q_RNIBG9H2_1_LC_5_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNIBG9H2_1_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNIBG9H2_1_LC_5_13_4 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNIBG9H2_1_LC_5_13_4  (
            .in0(N__11830),
            .in1(N__11651),
            .in2(N__11627),
            .in3(N__12728),
            .lcout(),
            .ltout(\Lab_UT.scdp.u1.N_539_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNIKMQ34_1_LC_5_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNIKMQ34_1_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNIKMQ34_1_LC_5_13_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNIKMQ34_1_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11586),
            .in3(N__11574),
            .lcout(),
            .ltout(\Lab_UT.scdp.N_426_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNI47LGA_1_LC_5_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNI47LGA_1_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNI47LGA_1_LC_5_13_6 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \Lab_UT.scdp.u0.q_RNI47LGA_1_LC_5_13_6  (
            .in0(N__12090),
            .in1(N__11544),
            .in2(N__11517),
            .in3(N__11775),
            .lcout(\Lab_UT.scdp.q_RNI47LGA_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_27_LC_5_13_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_27_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_27_LC_5_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_27_LC_5_13_7  (
            .in0(N__17931),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21078),
            .ce(N__12789),
            .sr(N__20851));
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_0_a2_0_x2_0_0_0_LC_5_14_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_0_a2_0_x2_0_0_0_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.b2a0.asciiHex_2_0_a2_0_x2_0_0_0_LC_5_14_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.b2a0.asciiHex_2_0_a2_0_x2_0_0_0_LC_5_14_0  (
            .in0(N__12807),
            .in1(N__11805),
            .in2(N__11886),
            .in3(N__12861),
            .lcout(\Lab_UT.scdp.b2a0.N_258_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIK3K3_1_LC_5_14_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIK3K3_1_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIK3K3_1_LC_5_14_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIK3K3_1_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__12798),
            .in2(_gnd_net_),
            .in3(N__11853),
            .lcout(\Lab_UT.scdp.d2eData_3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIMSEN_20_LC_5_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIMSEN_20_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIMSEN_20_LC_5_14_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIMSEN_20_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__12837),
            .in2(_gnd_net_),
            .in3(N__12543),
            .lcout(\Lab_UT.scdp.d2eData_3_0_a2_0_4 ),
            .ltout(\Lab_UT.scdp.d2eData_3_0_a2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI0Q781_4_LC_5_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI0Q781_4_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI0Q781_4_LC_5_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI0Q781_4_LC_5_14_6  (
            .in0(N__12806),
            .in1(N__12860),
            .in2(N__11799),
            .in3(N__17310),
            .lcout(\Lab_UT.scdp.N_246_i ),
            .ltout(\Lab_UT.scdp.N_246_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNI9Q034_1_LC_5_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNI9Q034_1_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNI9Q034_1_LC_5_14_7 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \Lab_UT.scdp.u0.q_RNI9Q034_1_LC_5_14_7  (
            .in0(N__12036),
            .in1(N__11769),
            .in2(N__11778),
            .in3(N__11972),
            .lcout(\Lab_UT.scdp.u0.L4_tx_data_0_a2_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNI41HI1_2_LC_5_15_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNI41HI1_2_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNI41HI1_2_LC_5_15_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.scdp.u1.q_RNI41HI1_2_LC_5_15_0  (
            .in0(N__12666),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12616),
            .lcout(\Lab_UT.scdp.N_256_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_2_LC_5_15_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_2_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_2_LC_5_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_2_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11763),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21072),
            .ce(N__12785),
            .sr(N__20853));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_10_LC_5_15_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_10_LC_5_15_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_10_LC_5_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_10_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14058),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21072),
            .ce(N__12785),
            .sr(N__20853));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIO7U41_2_LC_5_15_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIO7U41_2_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIO7U41_2_LC_5_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNIO7U41_2_LC_5_15_5  (
            .in0(N__12885),
            .in1(N__12105),
            .in2(N__12816),
            .in3(N__12099),
            .lcout(\Lab_UT.scdp.d2eData_3_2 ),
            .ltout(\Lab_UT.scdp.d2eData_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNI1L1F2_2_LC_5_15_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNI1L1F2_2_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNI1L1F2_2_LC_5_15_6 .LUT_INIT=16'b1010010111111111;
    LogicCell40 \Lab_UT.scdp.u1.q_RNI1L1F2_2_LC_5_15_6  (
            .in0(N__12667),
            .in1(_gnd_net_),
            .in2(N__12093),
            .in3(N__12081),
            .lcout(),
            .ltout(\Lab_UT.scdp.g0_0_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_RNIGMI45_1_LC_5_15_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_RNIGMI45_1_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_RNIGMI45_1_LC_5_15_7 .LUT_INIT=16'b1111001011110001;
    LogicCell40 \Lab_UT.scdp.u0.q_RNIGMI45_1_LC_5_15_7  (
            .in0(N__12047),
            .in1(N__11988),
            .in2(N__11979),
            .in3(N__11973),
            .lcout(\Lab_UT.scdp.g0_0_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_2_LC_6_3_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_2_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_2_LC_6_3_4 .LUT_INIT=16'b1100000001000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_2_LC_6_3_4  (
            .in0(N__19131),
            .in1(N__15457),
            .in2(N__11901),
            .in3(N__23209),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g1_1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_0_LC_6_3_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_0_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_0_LC_6_3_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_0_LC_6_3_5  (
            .in0(N__19493),
            .in1(N__23524),
            .in2(N__11910),
            .in3(N__12375),
            .lcout(\Lab_UT.scctrl.g1_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_6_0_LC_6_4_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_6_0_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_6_0_LC_6_4_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_6_0_LC_6_4_1  (
            .in0(N__16151),
            .in1(N__11907),
            .in2(N__14661),
            .in3(N__22968),
            .lcout(\Lab_UT.scctrl.N_399_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_o2_9_LC_6_4_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_o2_9_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_o2_9_LC_6_4_2 .LUT_INIT=16'b1110111011111011;
    LogicCell40 \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_o2_9_LC_6_4_2  (
            .in0(N__12165),
            .in1(N__14510),
            .in2(N__12188),
            .in3(N__18779),
            .lcout(\Lab_UT.scctrl.N_266i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_5_LC_6_4_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_5_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_5_LC_6_4_3 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_5_LC_6_4_3  (
            .in0(N__12891),
            .in1(N__19728),
            .in2(N__14660),
            .in3(N__22967),
            .lcout(\Lab_UT.scctrl.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_10_LC_6_4_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_10_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_10_LC_6_4_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_10_LC_6_4_4  (
            .in0(N__22966),
            .in1(N__18038),
            .in2(_gnd_net_),
            .in3(N__22041),
            .lcout(\Lab_UT.scctrl.N_319_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_5_LC_6_5_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_5_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_5_LC_6_5_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_5_LC_6_5_0  (
            .in0(N__21370),
            .in1(N__14766),
            .in2(N__12141),
            .in3(N__22286),
            .lcout(\Lab_UT.scctrl.N_414_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIVJ4S_LC_6_5_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIVJ4S_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIVJ4S_LC_6_5_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNIVJ4S_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__20585),
            .in2(_gnd_net_),
            .in3(N__21369),
            .lcout(\Lab_UT.scctrl.next_state_1_sqmuxa_10_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.state_1_ret_rep1_LC_6_5_2 .C_ON=1'b0;
    defparam \resetGen.state_1_ret_rep1_LC_6_5_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.state_1_ret_rep1_LC_6_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \resetGen.state_1_ret_rep1_LC_6_5_2  (
            .in0(N__22581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rst_i_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21113),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_0_LC_6_5_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_0_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_0_LC_6_5_4 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_RNIJFLD2_0_LC_6_5_4  (
            .in0(N__22042),
            .in1(N__19725),
            .in2(N__22464),
            .in3(N__22285),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_415_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNII8KJ5_3_LC_6_5_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNII8KJ5_3_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNII8KJ5_3_LC_6_5_5 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \Lab_UT.scctrl.state_2_RNII8KJ5_3_LC_6_5_5  (
            .in0(N__12117),
            .in1(N__23191),
            .in2(N__12120),
            .in3(N__22969),
            .lcout(\Lab_UT.scctrl.g1_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep2_RNITVAN_LC_6_5_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep2_RNITVAN_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep2_RNITVAN_LC_6_5_6 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep2_RNITVAN_LC_6_5_6  (
            .in0(N__22791),
            .in1(N__14652),
            .in2(N__18086),
            .in3(N__15443),
            .lcout(\Lab_UT.scctrl.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIIHUU_LC_6_5_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIIHUU_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIIHUU_LC_6_5_7 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNIIHUU_LC_6_5_7  (
            .in0(N__18905),
            .in1(N__22790),
            .in2(N__16316),
            .in3(N__18756),
            .lcout(\Lab_UT.scctrl.g0_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_2_LC_6_6_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_2_LC_6_6_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.shifter_ret_2_LC_6_6_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_2_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__13030),
            .in2(_gnd_net_),
            .in3(N__18782),
            .lcout(\Lab_UT.scctrl.N_241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21106),
            .ce(N__13447),
            .sr(N__20844));
    defparam \Lab_UT.scctrl.shifter_ret_14_LC_6_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_14_LC_6_6_1 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.scctrl.shifter_ret_14_LC_6_6_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_14_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__12111),
            .in2(_gnd_net_),
            .in3(N__14520),
            .lcout(\Lab_UT.scctrl.N_263_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21106),
            .ce(N__13447),
            .sr(N__20844));
    defparam \buart.Z_rx.shifter_ret_1_LC_6_6_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_1_LC_6_6_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_1_LC_6_6_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \buart.Z_rx.shifter_ret_1_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__17212),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21106),
            .ce(N__13447),
            .sr(N__20844));
    defparam \Lab_UT.scctrl.shifter_ret_5_LC_6_6_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_5_LC_6_6_3 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.scctrl.shifter_ret_5_LC_6_6_3 .LUT_INIT=16'b1111111011011101;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_5_LC_6_6_3  (
            .in0(N__18783),
            .in1(N__12164),
            .in2(N__12192),
            .in3(N__14521),
            .lcout(\Lab_UT.scctrl.N_266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21106),
            .ce(N__13447),
            .sr(N__20844));
    defparam \buart.Z_rx.shifter_ret_0_rep1_LC_6_6_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_0_rep1_LC_6_6_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_0_rep1_LC_6_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_0_rep1_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15083),
            .lcout(bu_rx_data_i_2_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21106),
            .ce(N__13447),
            .sr(N__20844));
    defparam \buart.Z_rx.shifter_0_4_LC_6_6_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_4_LC_6_6_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_4_LC_6_6_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_4_LC_6_6_5  (
            .in0(N__18784),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21106),
            .ce(N__13447),
            .sr(N__20844));
    defparam \Lab_UT.scdp.a2b.shifter_ret_RNISON11_LC_6_7_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.shifter_ret_RNISON11_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.shifter_ret_RNISON11_LC_6_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scdp.a2b.shifter_ret_RNISON11_LC_6_7_0  (
            .in0(N__13747),
            .in1(N__15181),
            .in2(N__12924),
            .in3(N__15071),
            .lcout(\Lab_UT.scdp.a2b.val_0_tz_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.a2b.val_i_o2_0_LC_6_7_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_i_o2_0_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_i_o2_0_LC_6_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scdp.a2b.val_i_o2_0_LC_6_7_1  (
            .in0(N__15072),
            .in1(N__13748),
            .in2(N__13517),
            .in3(N__15182),
            .lcout(\Lab_UT.scdp.a2b.N_280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_2_3_LC_6_7_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_3_LC_6_7_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_3_LC_6_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_3_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15074),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21099),
            .ce(N__13444),
            .sr(N__20839));
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_a2_3_LC_6_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_a2_3_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_a2_3_LC_6_7_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_a2_3_LC_6_7_4  (
            .in0(N__17129),
            .in1(N__13494),
            .in2(_gnd_net_),
            .in3(N__12150),
            .lcout(\Lab_UT.scctrl.N_472_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_4_LC_6_7_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_4_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_4_LC_6_7_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_4_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__12984),
            .in2(_gnd_net_),
            .in3(N__18788),
            .lcout(\Lab_UT.scctrl.N_241_reti ),
            .ltout(\Lab_UT.scctrl.N_241_reti_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_3_LC_6_7_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_LC_6_7_6 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.scctrl.shifter_ret_3_LC_6_7_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12144),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scctrl.N_241_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21099),
            .ce(N__13444),
            .sr(N__20839));
    defparam \buart.Z_rx.shifter_ret_0_LC_6_7_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_0_LC_6_7_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_0_LC_6_7_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_0_LC_6_7_7  (
            .in0(N__15073),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21099),
            .ce(N__13444),
            .sr(N__20839));
    defparam \Lab_UT.scctrl.shifter_ret_12_LC_6_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_12_LC_6_8_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.shifter_ret_12_LC_6_8_0 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_12_LC_6_8_0  (
            .in0(N__14937),
            .in1(N__17743),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scctrl.N_233_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21094),
            .ce(N__13443),
            .sr(N__20832));
    defparam \Lab_UT.scctrl.shifter_ret_12_RNIE3JF_LC_6_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_12_RNIE3JF_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_12_RNIE3JF_LC_6_8_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_12_RNIE3JF_LC_6_8_1  (
            .in0(N__12216),
            .in1(N__13404),
            .in2(_gnd_net_),
            .in3(N__12207),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_3_sqmuxa_i_0_i_o2_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNI0FVE3_LC_6_8_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNI0FVE3_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNI0FVE3_LC_6_8_2 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNI0FVE3_LC_6_8_2  (
            .in0(N__18904),
            .in1(N__12201),
            .in2(N__12195),
            .in3(N__14338),
            .lcout(\Lab_UT.scctrl.N_351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_8_LC_6_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_8_LC_6_8_3 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.scctrl.shifter_ret_8_LC_6_8_3 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_8_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17748),
            .in3(N__14936),
            .lcout(\Lab_UT.N_252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21094),
            .ce(N__13443),
            .sr(N__20832));
    defparam \buart.Z_rx.shifter_ret_3_LC_6_8_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_3_LC_6_8_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_3_LC_6_8_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_3_LC_6_8_4  (
            .in0(N__14938),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21094),
            .ce(N__13443),
            .sr(N__20832));
    defparam \buart.Z_rx.shifter_1_7_LC_6_8_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_7_LC_6_8_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_7_LC_6_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_1_7_LC_6_8_5  (
            .in0(N__17747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21094),
            .ce(N__13443),
            .sr(N__20832));
    defparam \buart.Z_rx.shifter_2_fast_6_LC_6_8_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_fast_6_LC_6_8_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_fast_6_LC_6_8_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_2_fast_6_LC_6_8_6  (
            .in0(N__14470),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buart__rx_shifter_2_fast_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21094),
            .ce(N__13443),
            .sr(N__20832));
    defparam \buart.Z_rx.shifter_ret_5_LC_6_8_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_5_LC_6_8_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_5_LC_6_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_5_LC_6_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14469),
            .lcout(bu_rx_data_i_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21094),
            .ce(N__13443),
            .sr(N__20832));
    defparam \buart.Z_rx.bitcount_es_1_LC_6_9_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_1_LC_6_9_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_1_LC_6_9_0 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_1_LC_6_9_0  (
            .in0(N__17694),
            .in1(N__13888),
            .in2(N__12240),
            .in3(N__13677),
            .lcout(buart__rx_bitcount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21089),
            .ce(N__12429),
            .sr(N__20840));
    defparam \buart.Z_rx.bitcount_es_2_LC_6_9_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_2_LC_6_9_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_2_LC_6_9_1 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_2_LC_6_9_1  (
            .in0(N__13889),
            .in1(N__17697),
            .in2(N__12228),
            .in3(N__13794),
            .lcout(\buart.Z_rx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21089),
            .ce(N__12429),
            .sr(N__20840));
    defparam CONSTANT_ONE_LUT4_LC_6_9_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_9_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_9_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(CONSTANT_ONE_NET_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_0_LC_6_9_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_0_LC_6_9_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_0_LC_6_9_3 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_0_LC_6_9_3  (
            .in0(N__13887),
            .in1(N__17696),
            .in2(N__12360),
            .in3(N__13865),
            .lcout(\buart.Z_rx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21089),
            .ce(N__12429),
            .sr(N__20840));
    defparam \buart.Z_rx.bitcount_es_3_LC_6_9_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_3_LC_6_9_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_3_LC_6_9_4 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_3_LC_6_9_4  (
            .in0(N__17695),
            .in1(N__13890),
            .in2(N__13827),
            .in3(N__12441),
            .lcout(\buart.Z_rx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21089),
            .ce(N__12429),
            .sr(N__20840));
    defparam \ufifo.emitcrlf_fsm.cstate_RNIQ8IQ3_0_LC_6_9_5 .C_ON=1'b0;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIQ8IQ3_0_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \ufifo.emitcrlf_fsm.cstate_RNIQ8IQ3_0_LC_6_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ufifo.emitcrlf_fsm.cstate_RNIQ8IQ3_0_LC_6_9_5  (
            .in0(N__12357),
            .in1(N__12345),
            .in2(_gnd_net_),
            .in3(N__12330),
            .lcout(utb_txdata_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_10_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__13861),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_10_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__13676),
            .in2(_gnd_net_),
            .in3(N__12231),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_10_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__13793),
            .in2(_gnd_net_),
            .in3(N__12219),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_10_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__13822),
            .in2(_gnd_net_),
            .in3(N__12435),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_4_LC_6_10_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_4_LC_6_10_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_4_LC_6_10_4 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_4_LC_6_10_4  (
            .in0(N__13886),
            .in1(N__17675),
            .in2(N__13731),
            .in3(N__12432),
            .lcout(buart__rx_bitcount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21083),
            .ce(N__12425),
            .sr(N__20843));
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIRA8MC_LC_6_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIRA8MC_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIRA8MC_LC_6_11_0 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_RNIRA8MC_LC_6_11_0  (
            .in0(N__12389),
            .in1(N__12399),
            .in2(N__15219),
            .in3(N__16736),
            .lcout(\Lab_UT.scctrl.next_state_rst_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_1_LC_6_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_1_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_1_LC_6_11_1 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_1_LC_6_11_1  (
            .in0(N__22187),
            .in1(N__22424),
            .in2(N__22059),
            .in3(N__22827),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_418_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI91NK6_0_2_LC_6_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI91NK6_0_2_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI91NK6_0_2_LC_6_11_2 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI91NK6_0_2_LC_6_11_2  (
            .in0(N__16703),
            .in1(N__19151),
            .in2(N__12402),
            .in3(N__23197),
            .lcout(\Lab_UT.scctrl.g0_2 ),
            .ltout(\Lab_UT.scctrl.g0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_3_LC_6_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_3_LC_6_11_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.next_state_3_LC_6_11_3 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \Lab_UT.scctrl.next_state_3_LC_6_11_3  (
            .in0(N__16737),
            .in1(N__15218),
            .in2(N__12393),
            .in3(N__12390),
            .lcout(\Lab_UT.scctrl.next_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21079),
            .ce(N__20900),
            .sr(N__20849));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_7_LC_6_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_7_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_7_LC_6_11_4 .LUT_INIT=16'b1010101010100010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_7_LC_6_11_4  (
            .in0(N__22828),
            .in1(N__22050),
            .in2(N__22454),
            .in3(N__22186),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_418_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_3_LC_6_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_3_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_3_LC_6_11_5 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_3_LC_6_11_5  (
            .in0(N__22188),
            .in1(N__14292),
            .in2(N__12378),
            .in3(N__21514),
            .lcout(\Lab_UT.scctrl.g1_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI6V451_2_LC_6_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI6V451_2_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI6V451_2_LC_6_11_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI6V451_2_LC_6_11_6  (
            .in0(N__22829),
            .in1(N__19152),
            .in2(N__21417),
            .in3(N__22051),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_39_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI6EDGH_2_LC_6_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI6EDGH_2_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI6EDGH_2_LC_6_11_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI6EDGH_2_LC_6_11_7  (
            .in0(N__12480),
            .in1(_gnd_net_),
            .in2(N__12363),
            .in3(N__15504),
            .lcout(\Lab_UT.state_1_RNI6EDGH_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_7_LC_6_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_7_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_7_LC_6_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_7_LC_6_12_0  (
            .in0(N__17043),
            .in1(N__17885),
            .in2(N__18395),
            .in3(N__16157),
            .lcout(\Lab_UT.scctrl.N_404_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNI9TOB1_LC_6_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNI9TOB1_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNI9TOB1_LC_6_12_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNI9TOB1_LC_6_12_1  (
            .in0(N__18356),
            .in1(N__20657),
            .in2(_gnd_net_),
            .in3(N__22052),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_22_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNI9C1NH_LC_6_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNI9C1NH_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNI9C1NH_LC_6_12_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNI9C1NH_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(N__15503),
            .in2(N__12531),
            .in3(N__12511),
            .lcout(\Lab_UT.state_1_ret_0_RNI9C1NH_0 ),
            .ltout(\Lab_UT.state_1_ret_0_RNI9C1NH_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.k3h.q_0_LC_6_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3h.q_0_LC_6_12_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3h.q_0_LC_6_12_3 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \Lab_UT.scdp.k3h.q_0_LC_6_12_3  (
            .in0(N__17617),
            .in1(N__12848),
            .in2(N__12528),
            .in3(N__18664),
            .lcout(\Lab_UT.scdp.key3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21076),
            .ce(),
            .sr(N__20820));
    defparam \Lab_UT.scdp.k3h.q_1_LC_6_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3h.q_1_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3h.q_1_LC_6_12_4 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \Lab_UT.scdp.k3h.q_1_LC_6_12_4  (
            .in0(N__17374),
            .in1(N__12524),
            .in2(N__18689),
            .in3(N__12512),
            .lcout(\Lab_UT.scdp.key3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21076),
            .ce(),
            .sr(N__20820));
    defparam \Lab_UT.scdp.k3h.q_2_LC_6_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3h.q_2_LC_6_12_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3h.q_2_LC_6_12_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.scdp.k3h.q_2_LC_6_12_5  (
            .in0(N__12513),
            .in1(N__18660),
            .in2(N__12497),
            .in3(N__16801),
            .lcout(\Lab_UT.scdp.key3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21076),
            .ce(),
            .sr(N__20820));
    defparam \Lab_UT.scdp.k0h.q_0_LC_6_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0h.q_0_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0h.q_0_LC_6_12_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k0h.q_0_LC_6_12_6  (
            .in0(N__18658),
            .in1(N__17616),
            .in2(N__12878),
            .in3(N__12476),
            .lcout(\Lab_UT.scdp.key0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21076),
            .ce(),
            .sr(N__20820));
    defparam \Lab_UT.scdp.k0h.q_1_LC_6_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0h.q_1_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0h.q_1_LC_6_12_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.scdp.k0h.q_1_LC_6_12_7  (
            .in0(N__12477),
            .in1(N__18659),
            .in2(N__12456),
            .in3(N__17375),
            .lcout(\Lab_UT.scdp.key0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21076),
            .ce(),
            .sr(N__20820));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_24_LC_6_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_24_LC_6_13_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_24_LC_6_13_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_24_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(N__16869),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21074),
            .ce(N__12787),
            .sr(N__20852));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_0_LC_6_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_0_LC_6_13_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_0_LC_6_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_0_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17577),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21074),
            .ce(N__12787),
            .sr(N__20852));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_16_LC_6_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_16_LC_6_13_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_16_LC_6_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_16_LC_6_13_3  (
            .in0(N__16908),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21074),
            .ce(N__12787),
            .sr(N__20852));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI9U1R_0_LC_6_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI9U1R_0_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI9U1R_0_LC_6_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_RNI9U1R_0_LC_6_13_4  (
            .in0(N__12759),
            .in1(N__12537),
            .in2(N__12753),
            .in3(N__12744),
            .lcout(\Lab_UT.scdp.d2eData_3_0 ),
            .ltout(\Lab_UT.scdp.d2eData_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNIJLK81_0_LC_6_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNIJLK81_0_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNIJLK81_0_LC_6_13_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNIJLK81_0_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12738),
            .in3(N__17262),
            .lcout(\Lab_UT.scdp.N_262_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNINM5R2_0_LC_6_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNINM5R2_0_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNINM5R2_0_LC_6_13_6 .LUT_INIT=16'b0000011001100000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNINM5R2_0_LC_6_13_6  (
            .in0(N__12626),
            .in1(N__12671),
            .in2(N__17268),
            .in3(N__12691),
            .lcout(\Lab_UT.scdp.u1.g0_0_i_a5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_RNINM5R2_0_0_LC_6_13_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_RNINM5R2_0_0_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u1.q_RNINM5R2_0_0_LC_6_13_7 .LUT_INIT=16'b0000011001100000;
    LogicCell40 \Lab_UT.scdp.u1.q_RNINM5R2_0_0_LC_6_13_7  (
            .in0(N__12690),
            .in1(N__17263),
            .in2(N__12672),
            .in3(N__12625),
            .lcout(\Lab_UT.scdp.u1.g0_0_i_a5_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_6_LC_6_14_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_6_LC_6_14_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_6_LC_6_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_6_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12591),
            .lcout(\Lab_UT.scdp.prng_lfsr_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21071),
            .ce(N__12786),
            .sr(N__20854));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_20_LC_6_14_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_20_LC_6_14_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_20_LC_6_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_20_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14087),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21071),
            .ce(N__12786),
            .sr(N__20854));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_8_LC_6_14_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_8_LC_6_14_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_8_LC_6_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_8_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14132),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21071),
            .ce(N__12786),
            .sr(N__20854));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_18_LC_6_14_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_18_LC_6_14_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_18_LC_6_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_18_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14072),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21071),
            .ce(N__12786),
            .sr(N__20854));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_4_LC_6_14_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_4_LC_6_14_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_4_LC_6_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_4_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12879),
            .lcout(\Lab_UT.scdp.prng_lfsr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21071),
            .ce(N__12786),
            .sr(N__20854));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_28_LC_6_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_28_LC_6_14_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_28_LC_6_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_28_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12852),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21071),
            .ce(N__12786),
            .sr(N__20854));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_11_LC_6_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_11_LC_6_14_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_11_LC_6_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_11_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14117),
            .lcout(\Lab_UT.scdp.prng_lfsr_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21071),
            .ce(N__12786),
            .sr(N__20854));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_26_LC_6_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_26_LC_6_14_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_26_LC_6_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_26_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16776),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21071),
            .ce(N__12786),
            .sr(N__20854));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_12_LC_6_15_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_12_LC_6_15_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_12_LC_6_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_12_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14018),
            .lcout(\Lab_UT.scdp.prng_lfsr_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21070),
            .ce(N__12784),
            .sr(N__20856));
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_9_LC_6_15_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_9_LC_6_15_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.lfsrInst.prng_lfsr_9_LC_6_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scdp.lfsrInst.prng_lfsr_9_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17334),
            .lcout(\Lab_UT.scdp.lfsrInst.prng_lfsrZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21070),
            .ce(N__12784),
            .sr(N__20856));
    defparam \Lab_UT.scctrl.sccEldByte_i_a2_0_LC_7_3_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.sccEldByte_i_a2_0_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.sccEldByte_i_a2_0_LC_7_3_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.sccEldByte_i_a2_0_LC_7_3_0  (
            .in0(N__12914),
            .in1(N__12897),
            .in2(N__13549),
            .in3(N__18803),
            .lcout(\Lab_UT.scctrl.N_385 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_a2_2_LC_7_3_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_a2_2_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_a2_2_LC_7_3_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.scctrl.next_state_1_sqmuxa_i_0_a2_2_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(N__18804),
            .in2(_gnd_net_),
            .in3(N__15106),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_534_reti_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_7_LC_7_3_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_7_LC_7_3_3 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.scctrl.shifter_ret_7_LC_7_3_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_7_LC_7_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13047),
            .in3(N__13044),
            .lcout(\Lab_UT.scctrl.N_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21137),
            .ce(N__13449),
            .sr(N__20855));
    defparam \Lab_UT.scdp.a2b.shifter_ret_LC_7_3_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.shifter_ret_LC_7_3_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scdp.a2b.shifter_ret_LC_7_3_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \Lab_UT.scdp.a2b.shifter_ret_LC_7_3_6  (
            .in0(_gnd_net_),
            .in1(N__17213),
            .in2(N__13550),
            .in3(N__13037),
            .lcout(\Lab_UT.N_540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21137),
            .ce(N__13449),
            .sr(N__20855));
    defparam \Lab_UT.scctrl.shifter_ret_13_LC_7_3_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_13_LC_7_3_7 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.scctrl.shifter_ret_13_LC_7_3_7 .LUT_INIT=16'b1011001110110011;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_13_LC_7_3_7  (
            .in0(N__15107),
            .in1(N__13537),
            .in2(N__17217),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scctrl.N_259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21137),
            .ce(N__13449),
            .sr(N__20855));
    defparam \Lab_UT.scctrl.state_1_RNO_8_0_LC_7_4_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_8_0_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_8_0_LC_7_4_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_8_0_LC_7_4_0  (
            .in0(N__16158),
            .in1(N__14514),
            .in2(_gnd_net_),
            .in3(N__13411),
            .lcout(\Lab_UT.scctrl.g0_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_2_0_LC_7_4_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_2_0_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_2_0_LC_7_4_1 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_2_0_LC_7_4_1  (
            .in0(N__12903),
            .in1(N__18245),
            .in2(N__18441),
            .in3(N__15455),
            .lcout(\Lab_UT.scctrl.g0_1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.sccEldByte_i_a2_0_1_LC_7_4_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.sccEldByte_i_a2_0_1_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.sccEldByte_i_a2_0_1_LC_7_4_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.scctrl.sccEldByte_i_a2_0_1_LC_7_4_2  (
            .in0(N__14926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15105),
            .lcout(\Lab_UT.scctrl.sccEldByte_i_a2_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_10_LC_7_4_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_10_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_10_LC_7_4_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_10_LC_7_4_3  (
            .in0(_gnd_net_),
            .in1(N__20577),
            .in2(_gnd_net_),
            .in3(N__21314),
            .lcout(\Lab_UT.scctrl.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_9_LC_7_4_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_9_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_9_LC_7_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_9_LC_7_4_4  (
            .in0(N__22034),
            .in1(N__18039),
            .in2(_gnd_net_),
            .in3(N__22975),
            .lcout(\Lab_UT.scctrl.N_319_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_1_LC_7_4_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_1_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_1_LC_7_4_6 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_1_LC_7_4_6  (
            .in0(N__13083),
            .in1(N__23706),
            .in2(N__23529),
            .in3(N__13065),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_1_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_LC_7_4_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_LC_7_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_ret_1_LC_7_4_7 .LUT_INIT=16'b0000010111111111;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_LC_7_4_7  (
            .in0(N__13104),
            .in1(_gnd_net_),
            .in2(N__13098),
            .in3(N__15456),
            .lcout(\Lab_UT.scctrl.N_235_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21129),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIUPHA1_LC_7_5_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIUPHA1_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIUPHA1_LC_7_5_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_RNIUPHA1_LC_7_5_0  (
            .in0(N__16576),
            .in1(N__13258),
            .in2(N__14939),
            .in3(N__14850),
            .lcout(\Lab_UT.scctrl.N_444_0 ),
            .ltout(\Lab_UT.scctrl.N_444_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_8_LC_7_5_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_8_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_8_LC_7_5_1 .LUT_INIT=16'b1111110011110010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_8_LC_7_5_1  (
            .in0(N__13355),
            .in1(N__15197),
            .in2(N__13095),
            .in3(N__15069),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_223_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_4_LC_7_5_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_4_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_4_LC_7_5_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_4_LC_7_5_2  (
            .in0(N__22268),
            .in1(N__13092),
            .in2(N__13086),
            .in3(N__21316),
            .lcout(\Lab_UT.scctrl.N_414_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.state_1_ret_fast_LC_7_5_3 .C_ON=1'b0;
    defparam \resetGen.state_1_ret_fast_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.state_1_ret_fast_LC_7_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \resetGen.state_1_ret_fast_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22580),
            .lcout(rst_i_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21124),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_4_LC_7_5_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_4_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_4_LC_7_5_4 .LUT_INIT=16'b1110110111101100;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNO_4_LC_7_5_4  (
            .in0(N__15070),
            .in1(N__13077),
            .in2(N__15201),
            .in3(N__13356),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_223_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_3_LC_7_5_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_3_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_3_LC_7_5_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNO_3_LC_7_5_5  (
            .in0(N__21317),
            .in1(N__18099),
            .in2(N__13071),
            .in3(N__22269),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_414_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_1_LC_7_5_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_1_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_1_LC_7_5_6 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNO_1_LC_7_5_6  (
            .in0(N__23696),
            .in1(N__23525),
            .in2(N__13068),
            .in3(N__13061),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_LC_7_5_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_ret_0_LC_7_5_7 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_LC_7_5_7  (
            .in0(N__15447),
            .in1(_gnd_net_),
            .in2(N__13050),
            .in3(N__15804),
            .lcout(\Lab_UT.scctrl.N_235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21124),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep1_RNIEMAA2_LC_7_6_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNIEMAA2_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNIEMAA2_LC_7_6_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep1_RNIEMAA2_LC_7_6_0  (
            .in0(N__16149),
            .in1(N__13116),
            .in2(N__20529),
            .in3(N__13128),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep1_RNIKQNN6_LC_7_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNIKQNN6_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNIKQNN6_LC_7_6_1 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep1_RNIKQNN6_LC_7_6_1  (
            .in0(N__23149),
            .in1(N__13953),
            .in2(N__13122),
            .in3(N__19316),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_0_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep2_RNI4KGMF_LC_7_6_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep2_RNI4KGMF_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep2_RNI4KGMF_LC_7_6_2 .LUT_INIT=16'b1111111110001111;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep2_RNI4KGMF_LC_7_6_2  (
            .in0(N__14653),
            .in1(N__14232),
            .in2(N__13119),
            .in3(N__19376),
            .lcout(\Lab_UT.scctrl.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNO_5_LC_7_6_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_5_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_5_LC_7_6_3 .LUT_INIT=16'b1000100000001000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNO_5_LC_7_6_3  (
            .in0(N__20528),
            .in1(N__16150),
            .in2(N__13200),
            .in3(N__22944),
            .lcout(\Lab_UT.scctrl.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI2SHF_LC_7_6_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI2SHF_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI2SHF_LC_7_6_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_2_RNI2SHF_LC_7_6_4  (
            .in0(N__13399),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16148),
            .lcout(\Lab_UT.scctrl.N_487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI8G3S_LC_7_6_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI8G3S_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI8G3S_LC_7_6_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_2_RNI8G3S_LC_7_6_5  (
            .in0(N__13250),
            .in1(N__13398),
            .in2(_gnd_net_),
            .in3(N__16988),
            .lcout(\Lab_UT.scctrl.N_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_15_LC_7_6_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_15_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_15_LC_7_6_6 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_15_LC_7_6_6  (
            .in0(N__16989),
            .in1(N__16147),
            .in2(N__13259),
            .in3(N__15878),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_2_0_0_a3_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_13_LC_7_6_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_13_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_13_LC_7_6_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_13_LC_7_6_7  (
            .in0(N__15952),
            .in1(N__14482),
            .in2(N__13110),
            .in3(N__14371),
            .lcout(\Lab_UT.scctrl.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_13_RNIORKJ_LC_7_7_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_13_RNIORKJ_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_13_RNIORKJ_LC_7_7_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_13_RNIORKJ_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__13219),
            .in2(_gnd_net_),
            .in3(N__21873),
            .lcout(\Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0 ),
            .ltout(\Lab_UT.scctrl.next_state_1_i_i_o2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep1_RNI5JDF1_LC_7_7_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNI5JDF1_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNI5JDF1_LC_7_7_1 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep1_RNI5JDF1_LC_7_7_1  (
            .in0(N__20521),
            .in1(N__19603),
            .in2(N__13107),
            .in3(N__16099),
            .lcout(\Lab_UT.scctrl.N_399 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI1JJ81_LC_7_7_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI1JJ81_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI1JJ81_LC_7_7_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_2_RNI1JJ81_LC_7_7_2  (
            .in0(N__16990),
            .in1(N__13254),
            .in2(N__19608),
            .in3(N__13400),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_i_o7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep2_RNIE3HB2_LC_7_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep2_RNIE3HB2_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep2_RNIE3HB2_LC_7_7_3 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep2_RNIE3HB2_LC_7_7_3  (
            .in0(N__14592),
            .in1(N__13272),
            .in2(N__13266),
            .in3(N__16100),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_12_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep2_RNIBDOL6_LC_7_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep2_RNIBDOL6_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep2_RNIBDOL6_LC_7_7_4 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep2_RNIBDOL6_LC_7_7_4  (
            .in0(N__13185),
            .in1(N__14208),
            .in2(N__13263),
            .in3(N__23128),
            .lcout(\Lab_UT.scctrl.g0_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNO_6_LC_7_7_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_6_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_6_LC_7_7_5 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNO_6_LC_7_7_5  (
            .in0(N__21875),
            .in1(N__13260),
            .in2(N__13224),
            .in3(N__16991),
            .lcout(\Lab_UT.scctrl.g0_1_i_a8_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIBUL06_LC_7_7_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIBUL06_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIBUL06_LC_7_7_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNIBUL06_LC_7_7_6  (
            .in0(N__21391),
            .in1(N__22250),
            .in2(N__20661),
            .in3(N__21479),
            .lcout(\Lab_UT.scctrl.N_401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNIQILS_0_LC_7_7_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNIQILS_0_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNIQILS_0_LC_7_7_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNIQILS_0_LC_7_7_7  (
            .in0(N__21874),
            .in1(N__19890),
            .in2(_gnd_net_),
            .in3(N__18265),
            .lcout(\Lab_UT.scctrl.N_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_9_LC_7_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_9_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_9_LC_7_8_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_9_LC_7_8_0  (
            .in0(N__15092),
            .in1(N__13179),
            .in2(_gnd_net_),
            .in3(N__15169),
            .lcout(\Lab_UT.scctrl.N_12_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_11_LC_7_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_11_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_11_LC_7_8_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_11_LC_7_8_1  (
            .in0(N__13173),
            .in1(N__13148),
            .in2(_gnd_net_),
            .in3(N__13563),
            .lcout(\Lab_UT.scctrl.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_0_RNI51T61_LC_7_8_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_0_RNI51T61_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_0_RNI51T61_LC_7_8_2 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_0_RNI51T61_LC_7_8_2  (
            .in0(N__13313),
            .in1(N__13172),
            .in2(N__13149),
            .in3(N__13562),
            .lcout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0 ),
            .ltout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_LC_7_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_LC_7_8_3 .LUT_INIT=16'b1111111110011000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_LC_7_8_3  (
            .in0(N__15168),
            .in1(N__15091),
            .in2(N__13359),
            .in3(N__13324),
            .lcout(\Lab_UT.scctrl.N_223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_1_LC_7_8_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_1_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_1_LC_7_8_4 .LUT_INIT=16'b1111101010101110;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_1_LC_7_8_4  (
            .in0(N__13325),
            .in1(N__13345),
            .in2(N__15120),
            .in3(N__15170),
            .lcout(\Lab_UT.scctrl.N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_0_LC_7_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_0_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_0_LC_7_8_5 .LUT_INIT=16'b1111111110011000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_RNIS5A43_0_LC_7_8_5  (
            .in0(N__15171),
            .in1(N__15096),
            .in2(N__13354),
            .in3(N__13326),
            .lcout(\Lab_UT.scctrl.N_223_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIESH11_LC_7_8_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIESH11_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIESH11_LC_7_8_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_RNIESH11_LC_7_8_6  (
            .in0(N__16241),
            .in1(N__14836),
            .in2(N__13314),
            .in3(N__13332),
            .lcout(\Lab_UT.scctrl.N_444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_ret_0_fast_LC_7_8_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_0_fast_LC_7_8_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_0_fast_LC_7_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_0_fast_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15097),
            .lcout(bu_rx_data_i_2_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21103),
            .ce(N__13445),
            .sr(N__20836));
    defparam \Lab_UT.scctrl.shifter_ret_LC_7_9_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_LC_7_9_0 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.scctrl.shifter_ret_LC_7_9_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__13290),
            .in2(_gnd_net_),
            .in3(N__13302),
            .lcout(\Lab_UT.scctrl.N_271_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21098),
            .ce(N__13442),
            .sr(N__20845));
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_5_LC_7_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_5_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_5_LC_7_9_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_5_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(N__13545),
            .in2(_gnd_net_),
            .in3(N__17196),
            .lcout(\Lab_UT.scctrl.N_219i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_RNI4H6R_LC_7_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_RNI4H6R_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_RNI4H6R_LC_7_9_2 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_RNI4H6R_LC_7_9_2  (
            .in0(N__13716),
            .in1(N__13670),
            .in2(N__13284),
            .in3(N__13412),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_1_sqmuxa_1_i_o2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_RNI7U912_LC_7_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_RNI7U912_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_RNI7U912_LC_7_9_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_RNI7U912_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13275),
            .in3(N__13764),
            .lcout(N_272),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_fast_0_LC_7_9_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_fast_0_LC_7_9_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_fast_0_LC_7_9_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_1_fast_0_LC_7_9_4  (
            .in0(N__17197),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buart__rx_shifter_1_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21098),
            .ce(N__13442),
            .sr(N__20845));
    defparam \buart.Z_rx.shifter_0_fast_2_LC_7_9_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_2_LC_7_9_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_2_LC_7_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_fast_2_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13547),
            .lcout(buart__rx_shifter_0_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21098),
            .ce(N__13442),
            .sr(N__20845));
    defparam \buart.Z_rx.shifter_ret_4_LC_7_9_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_4_LC_7_9_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_4_LC_7_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_4_LC_7_9_6  (
            .in0(N__13546),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21098),
            .ce(N__13442),
            .sr(N__20845));
    defparam \buart.Z_rx.shifter_1_0_LC_7_9_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_0_LC_7_9_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_0_LC_7_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_0_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17198),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21098),
            .ce(N__13442),
            .sr(N__20845));
    defparam \Lab_UT.scctrl.sccEldByte_i_o2_LC_7_10_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.sccEldByte_i_o2_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.sccEldByte_i_o2_LC_7_10_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \Lab_UT.scctrl.sccEldByte_i_o2_LC_7_10_0  (
            .in0(N__13673),
            .in1(N__14475),
            .in2(N__13730),
            .in3(N__13766),
            .lcout(\Lab_UT.scctrl.N_284 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_0_2_LC_7_10_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_0_2_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIPVCP_0_2_LC_7_10_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIPVCP_0_2_LC_7_10_1  (
            .in0(N__13791),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13820),
            .lcout(),
            .ltout(\buart.Z_rx.bitcountN11_15_i_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_0_LC_7_10_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_0_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_0_LC_7_10_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_0_0_LC_7_10_2  (
            .in0(N__13858),
            .in1(N__13726),
            .in2(N__13416),
            .in3(N__13675),
            .lcout(\buart.Z_rx.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI4KBA1_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI4KBA1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNI4KBA1_LC_7_10_3 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_2_RNI4KBA1_LC_7_10_3  (
            .in0(N__14474),
            .in1(N__13672),
            .in2(N__16146),
            .in3(N__13413),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_70_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_LC_7_10_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_LC_7_10_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_LC_7_10_4  (
            .in0(N__13721),
            .in1(N__13765),
            .in2(N__13362),
            .in3(N__15902),
            .lcout(\Lab_UT.scctrl.next_state_rst_0_3_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_4_LC_7_10_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_4_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_4_LC_7_10_5 .LUT_INIT=16'b0100111100001111;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOP0V3_4_LC_7_10_5  (
            .in0(N__13767),
            .in1(N__13722),
            .in2(N__17791),
            .in3(N__13674),
            .lcout(\buart.Z_rx.N_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNI3D361_2_LC_7_10_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNI3D361_2_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNI3D361_2_LC_7_10_6 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \buart.Z_rx.bitcount_es_RNI3D361_2_LC_7_10_6  (
            .in0(N__13857),
            .in1(_gnd_net_),
            .in2(N__13826),
            .in3(N__13790),
            .lcout(buart__rx_N_86_i_0_o2_1_0),
            .ltout(buart__rx_N_86_i_0_o2_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_8_RNIG4702_LC_7_10_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_8_RNIG4702_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_8_RNIG4702_LC_7_10_7 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_8_RNIG4702_LC_7_10_7  (
            .in0(N__13749),
            .in1(N__13717),
            .in2(N__13680),
            .in3(N__13671),
            .lcout(\Lab_UT.scctrl.N_261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.r4.q_0_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.r4.q_0_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.r4.q_0_LC_7_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scctrl.r4.q_0_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13610),
            .lcout(\Lab_UT.scctrl.r4.delay4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21087),
            .ce(),
            .sr(N__20821));
    defparam \Lab_UT.scctrl.r3.q_0_LC_7_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.r3.q_0_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.r3.q_0_LC_7_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scctrl.r3.q_0_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13590),
            .lcout(\Lab_UT.scctrl.delay3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21087),
            .ce(),
            .sr(N__20821));
    defparam \Lab_UT.scctrl.r1.q_0_LC_7_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.r1.q_0_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.r1.q_0_LC_7_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.scctrl.r1.q_0_LC_7_11_2  (
            .in0(N__15920),
            .in1(N__13584),
            .in2(N__21728),
            .in3(N__13578),
            .lcout(\Lab_UT.scctrl.delay1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21087),
            .ce(),
            .sr(N__20821));
    defparam \Lab_UT.scctrl.r2.q_0_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.r2.q_0_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.r2.q_0_LC_7_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scctrl.r2.q_0_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13596),
            .lcout(\Lab_UT.scctrl.delay2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21087),
            .ce(),
            .sr(N__20821));
    defparam \Lab_UT.scctrl.sccEldByte_i_a2_LC_7_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.sccEldByte_i_a2_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.sccEldByte_i_a2_LC_7_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.sccEldByte_i_a2_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__16138),
            .in2(_gnd_net_),
            .in3(N__15196),
            .lcout(\Lab_UT.scctrl.N_384 ),
            .ltout(\Lab_UT.scctrl.N_384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNIRGEB5_LC_7_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNIRGEB5_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNIRGEB5_LC_7_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNIRGEB5_LC_7_11_5  (
            .in0(N__13577),
            .in1(N__15919),
            .in2(N__13566),
            .in3(N__21717),
            .lcout(),
            .ltout(\Lab_UT.N_100_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u2.q_esr_ctle_7_LC_7_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u2.q_esr_ctle_7_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u2.q_esr_ctle_7_LC_7_11_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.scdp.u2.q_esr_ctle_7_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13908),
            .in3(N__20862),
            .lcout(\Lab_UT.scdp.u2.N_100_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_15_LC_7_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_15_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_15_LC_7_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_15_LC_7_12_0  (
            .in0(N__14633),
            .in1(N__17036),
            .in2(N__17896),
            .in3(N__16152),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_8_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_8_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_8_LC_7_12_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_8_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13896),
            .in3(N__19331),
            .lcout(\Lab_UT.scctrl.G_24_i_o7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_5_0_LC_7_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_5_0_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_5_0_LC_7_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_5_0_LC_7_12_2  (
            .in0(N__14634),
            .in1(N__17037),
            .in2(N__17894),
            .in3(N__16153),
            .lcout(\Lab_UT.scctrl.N_404_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_7_LC_7_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_7_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_7_LC_7_12_3 .LUT_INIT=16'b1010101010100010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_7_LC_7_12_3  (
            .in0(N__22819),
            .in1(N__22054),
            .in2(N__22462),
            .in3(N__22209),
            .lcout(\Lab_UT.scctrl.N_418_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_4_LC_7_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_4_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_4_LC_7_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNO_4_LC_7_12_4  (
            .in0(N__14636),
            .in1(N__17042),
            .in2(N__17895),
            .in3(N__16156),
            .lcout(\Lab_UT.scctrl.N_404_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_3_LC_7_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_3_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_3_LC_7_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_5_RNO_3_LC_7_12_5  (
            .in0(N__16154),
            .in1(N__17884),
            .in2(N__17053),
            .in3(N__14635),
            .lcout(\Lab_UT.scctrl.N_404_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_4_LC_7_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_4_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_4_LC_7_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNO_4_LC_7_12_6  (
            .in0(N__14637),
            .in1(N__17041),
            .in2(N__17897),
            .in3(N__16155),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_404_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_1_LC_7_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_1_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_1_LC_7_12_7 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNO_1_LC_7_12_7  (
            .in0(N__13944),
            .in1(N__19332),
            .in2(N__13893),
            .in3(N__21497),
            .lcout(\Lab_UT.scctrl.g0_2_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_3_RNI216C3_LC_7_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNI216C3_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNI216C3_LC_7_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_RNI216C3_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__15460),
            .in2(_gnd_net_),
            .in3(N__21495),
            .lcout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0 ),
            .ltout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_0_RNIIKTO3_LC_7_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_RNIIKTO3_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_0_RNIIKTO3_LC_7_13_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_RNIIKTO3_LC_7_13_1  (
            .in0(N__22046),
            .in1(_gnd_net_),
            .in2(N__14004),
            .in3(N__19729),
            .lcout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNI71T5A_LC_7_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNI71T5A_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNI71T5A_LC_7_13_2 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNI71T5A_LC_7_13_2  (
            .in0(N__15534),
            .in1(N__22199),
            .in2(N__14001),
            .in3(N__13968),
            .lcout(),
            .ltout(\Lab_UT.scctrl.un1_next_state_3_sqmuxa_2_0_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI0F8BG_0_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI0F8BG_0_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI0F8BG_0_LC_7_13_3 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI0F8BG_0_LC_7_13_3  (
            .in0(N__22201),
            .in1(N__21411),
            .in2(N__13962),
            .in3(N__13959),
            .lcout(\Lab_UT.scctrl.N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNIQILS_LC_7_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNIQILS_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNIQILS_LC_7_13_4 .LUT_INIT=16'b1111111100110000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNIQILS_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__22045),
            .in2(N__19906),
            .in3(N__18264),
            .lcout(\Lab_UT.scctrl.N_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_3_LC_7_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_3_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_3_LC_7_13_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNO_3_LC_7_13_5  (
            .in0(N__22200),
            .in1(N__20655),
            .in2(_gnd_net_),
            .in3(N__21410),
            .lcout(\Lab_UT.scctrl.g0_8_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_3_LC_7_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_3_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_3_LC_7_13_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNO_3_LC_7_13_6  (
            .in0(N__21412),
            .in1(N__20656),
            .in2(_gnd_net_),
            .in3(N__22202),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_1_LC_7_13_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_1_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_1_LC_7_13_7 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNO_1_LC_7_13_7  (
            .in0(N__21496),
            .in1(N__13938),
            .in2(N__13929),
            .in3(N__19333),
            .lcout(\Lab_UT.scctrl.g0_2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.k1h.q_2_LC_7_14_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1h.q_2_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1h.q_2_LC_7_14_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k1h.q_2_LC_7_14_0  (
            .in0(N__18665),
            .in1(N__16820),
            .in2(N__13925),
            .in3(N__17505),
            .lcout(\Lab_UT.scdp.key1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21075),
            .ce(),
            .sr(N__20824));
    defparam \Lab_UT.scdp.k1h.q_3_LC_7_14_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1h.q_3_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1h.q_3_LC_7_14_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.scdp.k1h.q_3_LC_7_14_1  (
            .in0(N__17506),
            .in1(N__18668),
            .in2(N__14150),
            .in3(N__18531),
            .lcout(\Lab_UT.scdp.key1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21075),
            .ce(),
            .sr(N__20824));
    defparam \Lab_UT.scdp.k1l.q_0_LC_7_14_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1l.q_0_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1l.q_0_LC_7_14_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k1l.q_0_LC_7_14_2  (
            .in0(N__18666),
            .in1(N__17626),
            .in2(N__14133),
            .in3(N__17354),
            .lcout(\Lab_UT.scdp.key1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21075),
            .ce(),
            .sr(N__20824));
    defparam \Lab_UT.scdp.k1l.q_3_LC_7_14_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1l.q_3_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1l.q_3_LC_7_14_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.scdp.k1l.q_3_LC_7_14_3  (
            .in0(N__17356),
            .in1(N__18669),
            .in2(N__14118),
            .in3(N__18532),
            .lcout(\Lab_UT.scdp.key1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21075),
            .ce(),
            .sr(N__20824));
    defparam \Lab_UT.scdp.k2h.q_2_LC_7_14_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2h.q_2_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2h.q_2_LC_7_14_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Lab_UT.scdp.k2h.q_2_LC_7_14_4  (
            .in0(N__18483),
            .in1(N__14099),
            .in2(N__18690),
            .in3(N__16824),
            .lcout(\Lab_UT.scdp.key2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21075),
            .ce(),
            .sr(N__20824));
    defparam \Lab_UT.scdp.k2h.q_0_LC_7_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2h.q_0_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2h.q_0_LC_7_14_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.scdp.k2h.q_0_LC_7_14_5  (
            .in0(N__17627),
            .in1(N__18670),
            .in2(N__14088),
            .in3(N__18482),
            .lcout(\Lab_UT.scdp.key2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21075),
            .ce(),
            .sr(N__20824));
    defparam \Lab_UT.scdp.k2l.q_2_LC_7_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2l.q_2_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2l.q_2_LC_7_14_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k2l.q_2_LC_7_14_6  (
            .in0(N__18667),
            .in1(N__16825),
            .in2(N__14073),
            .in3(N__17455),
            .lcout(\Lab_UT.scdp.key2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21075),
            .ce(),
            .sr(N__20824));
    defparam \Lab_UT.scdp.k1l.q_2_LC_7_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1l.q_2_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1l.q_2_LC_7_14_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \Lab_UT.scdp.k1l.q_2_LC_7_14_7  (
            .in0(N__17355),
            .in1(N__14051),
            .in2(N__16827),
            .in3(N__18674),
            .lcout(\Lab_UT.scdp.key1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21075),
            .ce(),
            .sr(N__20824));
    defparam \Lab_UT.scdp.k2h.q_1_LC_7_15_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2h.q_1_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2h.q_1_LC_7_15_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.scdp.k2h.q_1_LC_7_15_3  (
            .in0(N__18489),
            .in1(N__18688),
            .in2(N__14036),
            .in3(N__17402),
            .lcout(\Lab_UT.scdp.key2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21073),
            .ce(),
            .sr(N__20827));
    defparam \Lab_UT.scdp.k1h.q_0_LC_7_15_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1h.q_0_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1h.q_0_LC_7_15_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k1h.q_0_LC_7_15_5  (
            .in0(N__18687),
            .in1(N__17628),
            .in2(N__14019),
            .in3(N__17507),
            .lcout(\Lab_UT.scdp.key1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21073),
            .ce(),
            .sr(N__20827));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_16_LC_8_3_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_16_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_16_LC_8_3_2 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_16_LC_8_3_2  (
            .in0(N__20354),
            .in1(N__15747),
            .in2(_gnd_net_),
            .in3(N__16280),
            .lcout(\Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_8_LC_8_3_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_8_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_8_LC_8_3_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_8_LC_8_3_3  (
            .in0(N__14631),
            .in1(N__23453),
            .in2(N__18071),
            .in3(N__22804),
            .lcout(\Lab_UT.scctrl.N_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_3_0_LC_8_3_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_3_0_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_3_0_LC_8_3_4 .LUT_INIT=16'b0011001100010000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_3_0_LC_8_3_4  (
            .in0(N__18263),
            .in1(N__19392),
            .in2(N__14196),
            .in3(N__23190),
            .lcout(\Lab_UT.scctrl.g0_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep2_RNIN4FF_LC_8_3_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep2_RNIN4FF_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep2_RNIN4FF_LC_8_3_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep2_RNIN4FF_LC_8_3_5  (
            .in0(N__14630),
            .in1(N__18004),
            .in2(_gnd_net_),
            .in3(N__22803),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g1_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIVOU53_3_LC_8_3_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIVOU53_3_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIVOU53_3_LC_8_3_6 .LUT_INIT=16'b1000000010100000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIVOU53_3_LC_8_3_6  (
            .in0(N__15461),
            .in1(N__23189),
            .in2(N__14175),
            .in3(N__22971),
            .lcout(\Lab_UT.scctrl.g1_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_14_LC_8_4_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_14_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_14_LC_8_4_0 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_14_LC_8_4_0  (
            .in0(N__21305),
            .in1(N__16305),
            .in2(N__20605),
            .in3(N__14172),
            .lcout(\Lab_UT.scctrl.next_state_rst_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_0_LC_8_4_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_0_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_0_LC_8_4_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_0_LC_8_4_2  (
            .in0(N__14516),
            .in1(N__15896),
            .in2(N__15977),
            .in3(N__14384),
            .lcout(\Lab_UT.scctrl.N_290 ),
            .ltout(\Lab_UT.scctrl.N_290_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNO_2_LC_8_4_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_2_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_2_LC_8_4_3 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNO_2_LC_8_4_3  (
            .in0(N__18437),
            .in1(_gnd_net_),
            .in2(N__14166),
            .in3(N__18238),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNO_0_LC_8_4_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_0_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_0_LC_8_4_4 .LUT_INIT=16'b0010001000101110;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNO_0_LC_8_4_4  (
            .in0(N__20284),
            .in1(N__23496),
            .in2(N__14163),
            .in3(N__14259),
            .lcout(\Lab_UT.scctrl.next_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_4_0_LC_8_4_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_4_0_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_4_0_LC_8_4_5 .LUT_INIT=16'b0000000111111111;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_4_0_LC_8_4_5  (
            .in0(N__14385),
            .in1(N__14160),
            .in2(N__15903),
            .in3(N__18438),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_0_0_LC_8_4_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_0_0_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_0_0_LC_8_4_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_0_0_LC_8_4_6  (
            .in0(N__18702),
            .in1(N__14226),
            .in2(N__14220),
            .in3(N__14217),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_0_LC_8_4_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_0_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_0_LC_8_4_7 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.scctrl.state_1_0_LC_8_4_7  (
            .in0(N__23497),
            .in1(N__20285),
            .in2(N__14211),
            .in3(N__20183),
            .lcout(\Lab_UT.scctrl.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21138),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_1_LC_8_5_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_1_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_1_LC_8_5_0 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_RNIJFLD2_1_LC_8_5_0  (
            .in0(N__22031),
            .in1(N__19712),
            .in2(N__22420),
            .in3(N__22267),
            .lcout(\Lab_UT.scctrl.N_415_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNO_3_LC_8_5_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_3_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_3_LC_8_5_1 .LUT_INIT=16'b1011001100110011;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNO_3_LC_8_5_1  (
            .in0(N__18787),
            .in1(N__23572),
            .in2(N__18903),
            .in3(N__22700),
            .lcout(\Lab_UT.scctrl.g0_1_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNISO7C1_LC_8_5_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNISO7C1_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNISO7C1_LC_8_5_2 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNISO7C1_LC_8_5_2  (
            .in0(N__22698),
            .in1(N__18887),
            .in2(N__23589),
            .in3(N__18785),
            .lcout(\Lab_UT.scctrl.g0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_7_0_LC_8_5_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_7_0_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_7_0_LC_8_5_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_7_0_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__19847),
            .in2(_gnd_net_),
            .in3(N__22033),
            .lcout(\Lab_UT.scctrl.g3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep1_RNICQA1_LC_8_5_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNICQA1_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNICQA1_LC_8_5_4 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep1_RNICQA1_LC_8_5_4  (
            .in0(N__18203),
            .in1(N__20522),
            .in2(_gnd_net_),
            .in3(N__16306),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIBVSV_LC_8_5_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIBVSV_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIBVSV_LC_8_5_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNIBVSV_LC_8_5_5  (
            .in0(N__18786),
            .in1(N__18897),
            .in2(N__14184),
            .in3(N__22699),
            .lcout(\Lab_UT.scctrl.next_state_rst_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNO_4_LC_8_5_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_4_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_4_LC_8_5_6 .LUT_INIT=16'b0000000011011100;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNO_4_LC_8_5_6  (
            .in0(N__22032),
            .in1(N__18231),
            .in2(N__19873),
            .in3(N__23187),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_1_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNO_1_LC_8_5_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_1_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNO_1_LC_8_5_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNO_1_LC_8_5_7  (
            .in0(N__14181),
            .in1(N__14268),
            .in2(N__14262),
            .in3(N__19389),
            .lcout(\Lab_UT.scctrl.g0_1_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_12_LC_8_6_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_12_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_12_LC_8_6_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_12_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__19315),
            .in2(_gnd_net_),
            .in3(N__14253),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_24_i_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_6_LC_8_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_6_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_6_LC_8_6_1 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_6_LC_8_6_1  (
            .in0(N__18406),
            .in1(N__19369),
            .in2(N__14244),
            .in3(N__14241),
            .lcout(\Lab_UT.scctrl.G_24_i_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_11_LC_8_6_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_11_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_11_LC_8_6_2 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_11_LC_8_6_2  (
            .in0(N__20523),
            .in1(N__19577),
            .in2(_gnd_net_),
            .in3(N__19681),
            .lcout(\Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_6_LC_8_6_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_6_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_6_LC_8_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNO_6_LC_8_6_3  (
            .in0(N__14373),
            .in1(N__14518),
            .in2(N__15974),
            .in3(N__15892),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_290_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_2_LC_8_6_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_2_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_2_LC_8_6_4 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNO_2_LC_8_6_4  (
            .in0(N__18416),
            .in1(N__15695),
            .in2(N__14235),
            .in3(N__15543),
            .lcout(\Lab_UT.scctrl.g0_2_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_6_LC_8_6_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_6_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_6_LC_8_6_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNO_6_LC_8_6_5  (
            .in0(N__14374),
            .in1(N__14519),
            .in2(N__15975),
            .in3(N__15891),
            .lcout(\Lab_UT.scctrl.N_290_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_1_RNI4BLT2_0_LC_8_6_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_1_RNI4BLT2_0_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_1_RNI4BLT2_0_LC_8_6_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scctrl.state_ret_1_RNI4BLT2_0_LC_8_6_6  (
            .in0(N__14517),
            .in1(N__15879),
            .in2(N__18277),
            .in3(N__14372),
            .lcout(\Lab_UT.scctrl.N_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI6O741_2_LC_8_6_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI6O741_2_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI6O741_2_LC_8_6_7 .LUT_INIT=16'b1100110010001100;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI6O741_2_LC_8_6_7  (
            .in0(N__22741),
            .in1(N__15451),
            .in2(N__18433),
            .in3(N__19125),
            .lcout(\Lab_UT.scctrl.next_state_rst_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIECCO9_2_LC_8_7_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIECCO9_2_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIECCO9_2_LC_8_7_0 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIECCO9_2_LC_8_7_0  (
            .in0(N__19132),
            .in1(N__14550),
            .in2(N__14541),
            .in3(N__23150),
            .lcout(\Lab_UT.scctrl.next_state_rst_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_5_RNI1VIJ5_LC_8_7_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_5_RNI1VIJ5_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_5_RNI1VIJ5_LC_8_7_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_5_RNI1VIJ5_LC_8_7_1  (
            .in0(N__22284),
            .in1(N__16207),
            .in2(N__18058),
            .in3(N__21480),
            .lcout(\Lab_UT.scctrl.N_419_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep1_RNIHGED_LC_8_7_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNIHGED_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNIHGED_LC_8_7_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep1_RNIHGED_LC_8_7_2  (
            .in0(N__19573),
            .in1(N__20508),
            .in2(_gnd_net_),
            .in3(N__19687),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIDO8N1_LC_8_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIDO8N1_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIDO8N1_LC_8_7_3 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNIDO8N1_LC_8_7_3  (
            .in0(N__20643),
            .in1(N__23600),
            .in2(N__14544),
            .in3(N__21333),
            .lcout(\Lab_UT.scctrl.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_5_LC_8_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_5_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_5_LC_8_7_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_5_RNO_5_LC_8_7_4  (
            .in0(N__15901),
            .in1(N__14515),
            .in2(N__15976),
            .in3(N__14370),
            .lcout(\Lab_UT.scctrl.N_290_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_6_LC_8_7_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_6_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNO_6_LC_8_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNO_6_LC_8_7_5  (
            .in0(N__18028),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16206),
            .lcout(\Lab_UT.scctrl.g0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_fast_RNIKKMF_LC_8_7_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_fast_RNIKKMF_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_fast_RNIKKMF_LC_8_7_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_fast_RNIKKMF_LC_8_7_6  (
            .in0(N__19572),
            .in1(N__15743),
            .in2(_gnd_net_),
            .in3(N__20350),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_1_0_0_a2_2_0_0_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIGSGP1_LC_8_7_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIGSGP1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIGSGP1_LC_8_7_7 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNIGSGP1_LC_8_7_7  (
            .in0(N__20642),
            .in1(N__23599),
            .in2(N__14280),
            .in3(N__21332),
            .lcout(\Lab_UT.scctrl.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_LC_8_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_LC_8_8_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_13_LC_8_8_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_LC_8_8_0  (
            .in0(N__15663),
            .in1(N__14277),
            .in2(N__15624),
            .in3(N__20037),
            .lcout(\Lab_UT.N_245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21112),
            .ce(),
            .sr(N__20817));
    defparam \Lab_UT.scctrl.state_ret_12_LC_8_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_12_LC_8_8_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_12_LC_8_8_1 .LUT_INIT=16'b1110111110101011;
    LogicCell40 \Lab_UT.scctrl.state_ret_12_LC_8_8_1  (
            .in0(N__20038),
            .in1(N__23390),
            .in2(N__20287),
            .in3(N__14571),
            .lcout(\Lab_UT.scctrl.N_240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21112),
            .ce(),
            .sr(N__20817));
    defparam \Lab_UT.scctrl.state_ret_RNI3VN3G_LC_8_8_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_RNI3VN3G_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_RNI3VN3G_LC_8_8_2 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \Lab_UT.scctrl.state_ret_RNI3VN3G_LC_8_8_2  (
            .in0(N__15257),
            .in1(N__15312),
            .in2(N__18355),
            .in3(N__15287),
            .lcout(\Lab_UT.scctrl.next_state_rst ),
            .ltout(\Lab_UT.scctrl.next_state_rst_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_fast_LC_8_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_fast_LC_8_8_3 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_fast_LC_8_8_3 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \Lab_UT.scctrl.state_ret_fast_LC_8_8_3  (
            .in0(N__20268),
            .in1(_gnd_net_),
            .in2(N__14664),
            .in3(N__23392),
            .lcout(\Lab_UT.scctrl.state_i_1_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21112),
            .ce(),
            .sr(N__20817));
    defparam \Lab_UT.scctrl.state_ret_rep1_LC_8_8_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep1_LC_8_8_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_rep1_LC_8_8_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep1_LC_8_8_4  (
            .in0(N__23389),
            .in1(N__20269),
            .in2(_gnd_net_),
            .in3(N__16353),
            .lcout(\Lab_UT.scctrl.state_i_1_0_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21112),
            .ce(),
            .sr(N__20817));
    defparam \Lab_UT.scctrl.state_ret_5_LC_8_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_5_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_5_LC_8_8_5 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_5_LC_8_8_5  (
            .in0(N__20039),
            .in1(N__20276),
            .in2(N__16359),
            .in3(N__23391),
            .lcout(\Lab_UT.scctrl.N_240_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21112),
            .ce(),
            .sr(N__20817));
    defparam \Lab_UT.scctrl.state_ret_LC_8_8_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_LC_8_8_6 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_LC_8_8_6 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \Lab_UT.scctrl.state_ret_LC_8_8_6  (
            .in0(N__23388),
            .in1(N__20267),
            .in2(_gnd_net_),
            .in3(N__16352),
            .lcout(\Lab_UT.scctrl.state_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21112),
            .ce(),
            .sr(N__20817));
    defparam \Lab_UT.scctrl.state_ret_rep2_LC_8_8_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep2_LC_8_8_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_rep2_LC_8_8_7 .LUT_INIT=16'b0101010100001111;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep2_LC_8_8_7  (
            .in0(N__16354),
            .in1(_gnd_net_),
            .in2(N__20286),
            .in3(N__23393),
            .lcout(\Lab_UT.scctrl.state_i_1_0_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21112),
            .ce(),
            .sr(N__20817));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_0_LC_8_9_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_0_LC_8_9_0 .LUT_INIT=16'b0101001110101100;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_0_LC_8_9_0  (
            .in0(N__14805),
            .in1(N__19496),
            .in2(N__23452),
            .in3(N__20015),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_299_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_LC_8_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_4_LC_8_9_1 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_LC_8_9_1  (
            .in0(N__20184),
            .in1(N__15620),
            .in2(N__14574),
            .in3(N__14556),
            .lcout(Lab_UT_scctrl_N_223_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21104),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNI09OAV_0_LC_8_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNI09OAV_0_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNI09OAV_0_LC_8_9_2 .LUT_INIT=16'b1111111110001101;
    LogicCell40 \Lab_UT.scctrl.next_state_RNI09OAV_0_LC_8_9_2  (
            .in0(N__23352),
            .in1(N__14570),
            .in2(N__20283),
            .in3(N__20014),
            .lcout(\Lab_UT.scctrl.N_240_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_7_LC_8_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_7_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_7_LC_8_9_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_7_LC_8_9_3  (
            .in0(N__15792),
            .in1(N__15702),
            .in2(_gnd_net_),
            .in3(N__23351),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_2_0_0_a3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_3_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_3_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_3_LC_8_9_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_3_LC_8_9_4  (
            .in0(N__22842),
            .in1(N__14796),
            .in2(N__14715),
            .in3(N__14712),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_24_i_a3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_1_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_1_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_1_LC_8_9_5 .LUT_INIT=16'b1010101010111111;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_1_LC_8_9_5  (
            .in0(N__20016),
            .in1(N__14685),
            .in2(N__14703),
            .in3(N__14700),
            .lcout(\Lab_UT.scctrl.N_398i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_2_LC_8_9_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_2_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_2_LC_8_9_6 .LUT_INIT=16'b0101000000010000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_2_LC_8_9_6  (
            .in0(N__22841),
            .in1(N__14789),
            .in2(N__14694),
            .in3(N__22192),
            .lcout(\Lab_UT.scctrl.G_24_i_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_5_LC_8_9_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_5_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_5_LC_8_9_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_5_LC_8_9_7  (
            .in0(N__19495),
            .in1(N__20258),
            .in2(_gnd_net_),
            .in3(N__23350),
            .lcout(\Lab_UT.scctrl.G_24_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_4_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_4_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_4_LC_8_10_0 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_4_LC_8_10_0  (
            .in0(N__16365),
            .in1(N__14778),
            .in2(N__19008),
            .in3(N__14790),
            .lcout(\Lab_UT.scctrl.N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI9JP5A_1_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI9JP5A_1_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI9JP5A_1_LC_8_10_1 .LUT_INIT=16'b1111110010101000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI9JP5A_1_LC_8_10_1  (
            .in0(N__22189),
            .in1(N__22027),
            .in2(N__14676),
            .in3(N__14772),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIRHJAF_1_LC_8_10_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIRHJAF_1_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIRHJAF_1_LC_8_10_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIRHJAF_1_LC_8_10_2  (
            .in0(N__19434),
            .in1(N__23349),
            .in2(N__14667),
            .in3(N__16251),
            .lcout(\Lab_UT.scctrl.next_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_LC_8_10_3 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_RNIJFLD2_LC_8_10_3  (
            .in0(N__22191),
            .in1(N__22460),
            .in2(N__19730),
            .in3(N__22029),
            .lcout(\Lab_UT.scctrl.N_415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIBUL06_0_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIBUL06_0_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNIBUL06_0_LC_8_10_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNIBUL06_0_LC_8_10_4  (
            .in0(N__21501),
            .in1(N__21377),
            .in2(N__20662),
            .in3(N__22190),
            .lcout(\Lab_UT.scctrl.N_401_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_4_LC_8_10_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_4_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_4_LC_8_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_4_LC_8_10_5  (
            .in0(N__20651),
            .in1(N__22641),
            .in2(N__21409),
            .in3(N__21502),
            .lcout(\Lab_UT.scctrl.G_24_i_a7_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_8_LC_8_10_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_8_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_8_LC_8_10_6 .LUT_INIT=16'b1111111100100011;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_8_LC_8_10_6  (
            .in0(N__22028),
            .in1(N__18282),
            .in2(N__19945),
            .in3(N__23108),
            .lcout(\Lab_UT.scctrl.next_state_rst_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIN79O4_0_LC_8_10_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIN79O4_0_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIN79O4_0_LC_8_10_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIN79O4_0_LC_8_10_7  (
            .in0(N__23348),
            .in1(N__21390),
            .in2(N__18954),
            .in3(N__21500),
            .lcout(\Lab_UT.scctrl.G_15_0_a10_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_9_LC_8_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_9_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_9_LC_8_11_0 .LUT_INIT=16'b0111111100001111;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_9_LC_8_11_0  (
            .in0(N__21499),
            .in1(N__16212),
            .in2(N__19156),
            .in3(N__23117),
            .lcout(\Lab_UT.scctrl.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNIKFLC4_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNIKFLC4_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNIKFLC4_LC_8_11_1 .LUT_INIT=16'b0000011111111111;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNIKFLC4_LC_8_11_1  (
            .in0(N__21388),
            .in1(N__22037),
            .in2(N__19941),
            .in3(N__21498),
            .lcout(\Lab_UT.scctrl.g0_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNI4P8F2_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNI4P8F2_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNI4P8F2_LC_8_11_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.scctrl.state_1_2_rep1_RNI4P8F2_LC_8_11_2  (
            .in0(N__20451),
            .in1(N__16211),
            .in2(_gnd_net_),
            .in3(N__22175),
            .lcout(\Lab_UT.scctrl.g0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_3_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_3_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_3_LC_8_11_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_3_LC_8_11_3  (
            .in0(N__22177),
            .in1(N__14762),
            .in2(N__19157),
            .in3(N__16210),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_419_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_0_LC_8_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_0_LC_8_11_4 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_0_LC_8_11_4  (
            .in0(N__19492),
            .in1(N__23463),
            .in2(N__14745),
            .in3(N__15225),
            .lcout(\Lab_UT.scctrl.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_6_LC_8_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_6_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_6_LC_8_11_5 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_6_LC_8_11_5  (
            .in0(N__21389),
            .in1(N__20647),
            .in2(N__14730),
            .in3(N__15450),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_2_LC_8_11_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_2_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_2_RNO_2_LC_8_11_6 .LUT_INIT=16'b0101000000010000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_2_RNO_2_LC_8_11_6  (
            .in0(N__15234),
            .in1(N__19144),
            .in2(N__15228),
            .in3(N__23118),
            .lcout(\Lab_UT.scctrl.g0_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_0_LC_8_11_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_0_LC_8_11_7 .LUT_INIT=16'b1100100011001100;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_0_LC_8_11_7  (
            .in0(N__22176),
            .in1(N__22792),
            .in2(N__22461),
            .in3(N__22036),
            .lcout(\Lab_UT.scctrl.N_418_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_3_RNI7ARC1_LC_8_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNI7ARC1_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNI7ARC1_LC_8_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_RNI7ARC1_LC_8_12_0  (
            .in0(N__14852),
            .in1(N__16560),
            .in2(N__14949),
            .in3(N__17890),
            .lcout(\Lab_UT.scctrl.N_444_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_3_RNI7ARC1_0_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNI7ARC1_0_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNI7ARC1_0_LC_8_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_RNI7ARC1_0_LC_8_12_1  (
            .in0(N__14941),
            .in1(N__16559),
            .in2(N__17898),
            .in3(N__14851),
            .lcout(\Lab_UT.scctrl.N_444_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_7_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_7_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_7_LC_8_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_7_LC_8_12_2  (
            .in0(N__16208),
            .in1(N__15195),
            .in2(N__20456),
            .in3(N__15129),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_24_i_a6_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_3_LC_8_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_3_LC_8_12_3 .LUT_INIT=16'b1101110011011000;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_3_LC_8_12_3  (
            .in0(N__22236),
            .in1(N__22826),
            .in2(N__14964),
            .in3(N__15243),
            .lcout(\Lab_UT.scctrl.G_24_i_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_4_LC_8_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_4_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_4_LC_8_12_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_4_LC_8_12_4  (
            .in0(N__16209),
            .in1(N__17891),
            .in2(N__18087),
            .in3(N__22235),
            .lcout(\Lab_UT.scctrl.G_24_i_a6_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_5_LC_8_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_5_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_5_LC_8_12_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_5_LC_8_12_5  (
            .in0(N__16561),
            .in1(N__14961),
            .in2(N__14948),
            .in3(N__14853),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_1_LC_8_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_1_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_1_LC_8_12_6 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_1_LC_8_12_6  (
            .in0(N__14820),
            .in1(N__14814),
            .in2(N__14808),
            .in3(N__15318),
            .lcout(\Lab_UT.scctrl.next_state_rst_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_2_LC_8_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_2_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_2_LC_8_12_7 .LUT_INIT=16'b1101110111111101;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_2_LC_8_12_7  (
            .in0(N__23607),
            .in1(N__16029),
            .in2(N__18085),
            .in3(N__23119),
            .lcout(\Lab_UT.scctrl.G_24_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_0_LC_8_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_0_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.next_state_0_LC_8_13_0 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \Lab_UT.scctrl.next_state_0_LC_8_13_0  (
            .in0(N__15311),
            .in1(N__15291),
            .in2(N__18439),
            .in3(N__15264),
            .lcout(\Lab_UT.scctrl.next_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21081),
            .ce(N__20899),
            .sr(N__20857));
    defparam \Lab_UT.scctrl.state_ret_RNIKML91_LC_8_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_RNIKML91_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_RNIKML91_LC_8_13_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_RNIKML91_LC_8_13_1  (
            .in0(N__16013),
            .in1(N__18420),
            .in2(_gnd_net_),
            .in3(N__22057),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_170_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_RNIK5UKH_LC_8_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_RNIK5UKH_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_RNIK5UKH_LC_8_13_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.scctrl.state_ret_RNIK5UKH_LC_8_13_2  (
            .in0(N__15498),
            .in1(_gnd_net_),
            .in2(N__15246),
            .in3(N__17457),
            .lcout(\Lab_UT.state_ret_RNIK5UKH_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_12_RNIUVHQG_LC_8_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_12_RNIUVHQG_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_12_RNIUVHQG_LC_8_13_3 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_12_RNIUVHQG_LC_8_13_3  (
            .in0(N__17952),
            .in1(N__19814),
            .in2(N__16017),
            .in3(N__15499),
            .lcout(\Lab_UT.state_ret_12_RNIUVHQG_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_8_LC_8_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_8_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_8_LC_8_13_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_8_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__22442),
            .in2(_gnd_net_),
            .in3(N__22053),
            .lcout(\Lab_UT.scctrl.G_24_i_o6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_12_RNI2D6E_LC_8_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_12_RNI2D6E_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_12_RNI2D6E_LC_8_13_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.scctrl.state_ret_12_RNI2D6E_LC_8_13_5  (
            .in0(N__19813),
            .in1(N__19158),
            .in2(_gnd_net_),
            .in3(N__22802),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_17_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_12_RNI2SEPG_LC_8_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_12_RNI2SEPG_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_12_RNI2SEPG_LC_8_13_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.scctrl.state_ret_12_RNI2SEPG_LC_8_13_6  (
            .in0(N__15497),
            .in1(_gnd_net_),
            .in2(N__15237),
            .in3(N__17358),
            .lcout(\Lab_UT.state_ret_12_RNI2SEPG_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI2IGHH_0_LC_8_13_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI2IGHH_0_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI2IGHH_0_LC_8_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI2IGHH_0_LC_8_13_7  (
            .in0(N__18488),
            .in1(N__15990),
            .in2(_gnd_net_),
            .in3(N__15496),
            .lcout(\Lab_UT.state_1_RNI2IGHH_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIOII81_2_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIOII81_2_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIOII81_2_LC_8_14_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIOII81_2_LC_8_14_1  (
            .in0(N__19154),
            .in1(N__22823),
            .in2(N__18440),
            .in3(N__22055),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_20_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIO1RJH_2_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIO1RJH_2_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIO1RJH_2_LC_8_14_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIO1RJH_2_LC_8_14_2  (
            .in0(N__17549),
            .in1(_gnd_net_),
            .in2(N__15537),
            .in3(N__15494),
            .lcout(\Lab_UT.state_1_RNIO1RJH_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNILCGA1_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNILCGA1_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNILCGA1_LC_8_14_3 .LUT_INIT=16'b0001000111110001;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNILCGA1_LC_8_14_3  (
            .in0(N__19153),
            .in1(N__22822),
            .in2(N__20691),
            .in3(N__16012),
            .lcout(\Lab_UT.scctrl.N_277 ),
            .ltout(\Lab_UT.scctrl.N_277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIR2443_LC_8_14_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIR2443_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIR2443_LC_8_14_4 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNIR2443_LC_8_14_4  (
            .in0(N__22976),
            .in1(N__15510),
            .in2(N__15528),
            .in3(N__18906),
            .lcout(N_67),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_RNIVRBS_LC_8_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_RNIVRBS_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_RNIVRBS_LC_8_14_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_RNIVRBS_LC_8_14_5  (
            .in0(N__18427),
            .in1(N__22825),
            .in2(_gnd_net_),
            .in3(N__22056),
            .lcout(\Lab_UT.scctrl.N_355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNI2KLS_LC_8_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNI2KLS_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNI2KLS_LC_8_14_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNI2KLS_LC_8_14_6  (
            .in0(N__22824),
            .in1(N__20690),
            .in2(_gnd_net_),
            .in3(N__19155),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_27_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNI23U7H_LC_8_14_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNI23U7H_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNI23U7H_LC_8_14_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNI23U7H_LC_8_14_7  (
            .in0(N__15495),
            .in1(_gnd_net_),
            .in2(N__15465),
            .in3(N__17508),
            .lcout(\Lab_UT.state_1_ret_3_RNI23U7H_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_3_LC_9_3_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_3_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_3_LC_9_3_1 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_3_LC_9_3_1  (
            .in0(N__23488),
            .in1(N__15462),
            .in2(N__15327),
            .in3(N__19340),
            .lcout(\Lab_UT.scctrl.G_18_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_2_LC_9_4_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_2_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_2_LC_9_4_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.scctrl.state_1_2_LC_9_4_0  (
            .in0(N__15567),
            .in1(N__15588),
            .in2(N__23708),
            .in3(N__23494),
            .lcout(\Lab_UT.scctrl.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20826));
    defparam \Lab_UT.scctrl.state_1_fast_2_LC_9_4_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_fast_2_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_fast_2_LC_9_4_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Lab_UT.scctrl.state_1_fast_2_LC_9_4_1  (
            .in0(N__23491),
            .in1(N__23705),
            .in2(N__15597),
            .in3(N__15570),
            .lcout(\Lab_UT.scctrl.state_fast_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20826));
    defparam \Lab_UT.scctrl.state_1_2_rep1_LC_9_4_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_2_rep1_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_2_rep1_LC_9_4_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.scctrl.state_1_2_rep1_LC_9_4_2  (
            .in0(N__15568),
            .in1(N__15589),
            .in2(N__23709),
            .in3(N__23495),
            .lcout(\Lab_UT.scctrl.state_2_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20826));
    defparam \Lab_UT.scctrl.state_ret_0_RNI1ME69_LC_9_4_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_RNI1ME69_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_0_RNI1ME69_LC_9_4_3 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_RNI1ME69_LC_9_4_3  (
            .in0(N__22296),
            .in1(N__15654),
            .in2(N__15711),
            .in3(N__21522),
            .lcout(\Lab_UT.scctrl.g1_2_0 ),
            .ltout(\Lab_UT.scctrl.g1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNI3K1MC_2_LC_9_4_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNI3K1MC_2_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNI3K1MC_2_LC_9_4_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Lab_UT.scctrl.next_state_RNI3K1MC_2_LC_9_4_4  (
            .in0(N__23697),
            .in1(N__15587),
            .in2(N__15648),
            .in3(N__23489),
            .lcout(\Lab_UT.scctrl.next_stateZ0Z_2 ),
            .ltout(\Lab_UT.scctrl.next_stateZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_LC_9_4_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_LC_9_4_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_11_LC_9_4_5 .LUT_INIT=16'b0001111110111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_LC_9_4_5  (
            .in0(N__23492),
            .in1(N__19530),
            .in2(N__15645),
            .in3(N__15641),
            .lcout(\Lab_UT.scctrl.N_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20826));
    defparam \Lab_UT.scctrl.state_ret_1_LC_9_4_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_1_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_1_LC_9_4_6 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_1_LC_9_4_6  (
            .in0(N__15642),
            .in1(N__23493),
            .in2(N__19536),
            .in3(N__15613),
            .lcout(\Lab_UT.scctrl.N_296_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20826));
    defparam \Lab_UT.scctrl.state_1_2_rep2_LC_9_4_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_2_rep2_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_2_rep2_LC_9_4_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Lab_UT.scctrl.state_1_2_rep2_LC_9_4_7  (
            .in0(N__23490),
            .in1(N__23704),
            .in2(N__15596),
            .in3(N__15569),
            .lcout(\Lab_UT.scctrl.state_2_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21143),
            .ce(),
            .sr(N__20826));
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_4_LC_9_5_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_4_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_4_LC_9_5_0 .LUT_INIT=16'b1111111100100011;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_5_RNO_4_LC_9_5_0  (
            .in0(N__21996),
            .in1(N__18230),
            .in2(N__19944),
            .in3(N__23186),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_2_LC_9_5_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_2_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_2_LC_9_5_1 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_5_RNO_2_LC_9_5_1  (
            .in0(N__18432),
            .in1(N__15698),
            .in2(N__15555),
            .in3(N__15552),
            .lcout(\Lab_UT.scctrl.g0_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_5_LC_9_5_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_5_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_5_LC_9_5_2 .LUT_INIT=16'b1111111100100011;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNO_5_LC_9_5_2  (
            .in0(N__21993),
            .in1(N__18225),
            .in2(N__19942),
            .in3(N__23183),
            .lcout(\Lab_UT.scctrl.next_state_rst_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_5_LC_9_5_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_5_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_5_LC_9_5_3 .LUT_INIT=16'b1010111110101011;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNO_5_LC_9_5_3  (
            .in0(N__23185),
            .in1(N__19926),
            .in2(N__18259),
            .in3(N__21997),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_4_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_2_LC_9_5_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_2_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_2_LC_9_5_4 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNO_2_LC_9_5_4  (
            .in0(N__15697),
            .in1(N__18431),
            .in2(N__15720),
            .in3(N__15717),
            .lcout(\Lab_UT.scctrl.g0_2_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_2_rep2_RNI2S7K1_LC_9_5_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_2_rep2_RNI2S7K1_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_2_rep2_RNI2S7K1_LC_9_5_5 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \Lab_UT.scctrl.state_1_2_rep2_RNI2S7K1_LC_9_5_5  (
            .in0(N__21315),
            .in1(N__21994),
            .in2(N__18054),
            .in3(N__22918),
            .lcout(\Lab_UT.scctrl.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNI1HVT2_LC_9_5_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNI1HVT2_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNI1HVT2_LC_9_5_6 .LUT_INIT=16'b1111111100100011;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNI1HVT2_LC_9_5_6  (
            .in0(N__21995),
            .in1(N__18226),
            .in2(N__19943),
            .in3(N__23184),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_RNI227Q7_LC_9_5_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_RNI227Q7_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_RNI227Q7_LC_9_5_7 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_RNI227Q7_LC_9_5_7  (
            .in0(N__18430),
            .in1(N__15696),
            .in2(N__15672),
            .in3(N__15669),
            .lcout(\Lab_UT.scctrl.g0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIB2MFC_3_LC_9_6_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIB2MFC_3_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIB2MFC_3_LC_9_6_0 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIB2MFC_3_LC_9_6_0  (
            .in0(N__19242),
            .in1(N__19521),
            .in2(N__23498),
            .in3(N__15787),
            .lcout(\Lab_UT.scctrl.next_state_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_fast_3_LC_9_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_fast_3_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_2_fast_3_LC_9_6_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \Lab_UT.scctrl.state_2_fast_3_LC_9_6_1  (
            .in0(N__15790),
            .in1(N__23426),
            .in2(N__19535),
            .in3(N__19245),
            .lcout(\Lab_UT.scctrl.state_fast_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(),
            .sr(N__20823));
    defparam \Lab_UT.scctrl.state_2_3_rep1_LC_9_6_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_3_rep1_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_2_3_rep1_LC_9_6_2 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \Lab_UT.scctrl.state_2_3_rep1_LC_9_6_2  (
            .in0(N__19244),
            .in1(N__19525),
            .in2(N__23499),
            .in3(N__15789),
            .lcout(\Lab_UT.scctrl.state_3_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(),
            .sr(N__20823));
    defparam \Lab_UT.scctrl.state_2_3_LC_9_6_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_3_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_2_3_LC_9_6_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \Lab_UT.scctrl.state_2_3_LC_9_6_3  (
            .in0(N__15788),
            .in1(N__23425),
            .in2(N__19534),
            .in3(N__19243),
            .lcout(\Lab_UT.scctrl.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(),
            .sr(N__20823));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_2_LC_9_6_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_2_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_2_LC_9_6_4 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNO_2_LC_9_6_4  (
            .in0(N__22290),
            .in1(N__22400),
            .in2(N__22044),
            .in3(N__22737),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_418_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_0_LC_9_6_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_0_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_0_LC_9_6_5 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNO_0_LC_9_6_5  (
            .in0(N__19520),
            .in1(N__23421),
            .in2(N__15807),
            .in3(N__19241),
            .lcout(\Lab_UT.scctrl.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_6_LC_9_6_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_6_LC_9_6_6 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_6_LC_9_6_6 .LUT_INIT=16'b1111001101010011;
    LogicCell40 \Lab_UT.scctrl.state_ret_6_LC_9_6_6  (
            .in0(N__19246),
            .in1(N__19529),
            .in2(N__23500),
            .in3(N__15791),
            .lcout(\Lab_UT.scctrl.state_i_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21130),
            .ce(),
            .sr(N__20823));
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_LC_9_6_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_LC_9_6_7 .LUT_INIT=16'b1010101010100010;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_7_RNIPFLD2_LC_9_6_7  (
            .in0(N__22736),
            .in1(N__21989),
            .in2(N__22440),
            .in3(N__22289),
            .lcout(\Lab_UT.scctrl.N_418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_0_LC_9_7_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_LC_9_7_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_0_LC_9_7_0 .LUT_INIT=16'b1011000110111011;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_LC_9_7_0  (
            .in0(N__23433),
            .in1(N__23691),
            .in2(N__15765),
            .in3(N__18113),
            .lcout(\Lab_UT.scctrl.state_i_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21125),
            .ce(),
            .sr(N__20822));
    defparam \Lab_UT.scctrl.state_ret_0_fast_LC_9_7_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_fast_LC_9_7_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.scctrl.state_ret_0_fast_LC_9_7_1 .LUT_INIT=16'b1101110100001111;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_fast_LC_9_7_1  (
            .in0(N__18114),
            .in1(N__15764),
            .in2(N__23707),
            .in3(N__23434),
            .lcout(\Lab_UT.scctrl.state_ret_0_fastZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21125),
            .ce(),
            .sr(N__20822));
    defparam \Lab_UT.scctrl.state_ret_0_RNIKR11_LC_9_7_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_RNIKR11_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_0_RNIKR11_LC_9_7_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_RNIKR11_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__23394),
            .in2(_gnd_net_),
            .in3(N__19669),
            .lcout(\Lab_UT.scctrl.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_11_LC_9_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_11_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_11_LC_9_7_3 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_11_LC_9_7_3  (
            .in0(N__15742),
            .in1(_gnd_net_),
            .in2(N__23487),
            .in3(N__22769),
            .lcout(\Lab_UT.scctrl.G_18_i_a9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_10_LC_9_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_10_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_10_LC_9_7_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_10_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__16279),
            .in2(_gnd_net_),
            .in3(N__15741),
            .lcout(),
            .ltout(\Lab_UT.scctrl.state_ret_4_RNOZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNO_6_LC_9_7_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_6_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNO_6_LC_9_7_5 .LUT_INIT=16'b0011000111110101;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNO_6_LC_9_7_5  (
            .in0(N__20520),
            .in1(N__20641),
            .in2(N__16032),
            .in3(N__21364),
            .lcout(\Lab_UT.scctrl.state_ret_4_RNOZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_0_RNIJOQD_LC_9_7_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_RNIJOQD_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_0_RNIJOQD_LC_9_7_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_RNIJOQD_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__19670),
            .in2(_gnd_net_),
            .in3(N__22888),
            .lcout(\Lab_UT.scctrl.N_295 ),
            .ltout(\Lab_UT.scctrl.N_295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI23861_0_LC_9_7_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI23861_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI23861_0_LC_9_7_7 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI23861_0_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__21365),
            .in2(N__15993),
            .in3(N__21960),
            .lcout(\Lab_UT.scctrl.N_40_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_1_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_1_LC_9_8_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_2_RNID9MC3_1_LC_9_8_0  (
            .in0(N__15978),
            .in1(N__15924),
            .in2(_gnd_net_),
            .in3(N__15900),
            .lcout(\Lab_UT.scctrl.next_state_rst_0_3_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNIJJLN1_LC_9_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNIJJLN1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNIJJLN1_LC_9_8_1 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_2_rep1_RNIJJLN1_LC_9_8_1  (
            .in0(N__21974),
            .in1(N__20452),
            .in2(N__16575),
            .in3(N__16104),
            .lcout(\Lab_UT.scctrl.N_408 ),
            .ltout(\Lab_UT.scctrl.N_408_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_16_LC_9_8_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_16_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_16_LC_9_8_2 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_16_LC_9_8_2  (
            .in0(N__16040),
            .in1(N__16218),
            .in2(N__15837),
            .in3(N__23179),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_i_a8_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_9_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_9_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_9_LC_9_8_3 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_9_LC_9_8_3  (
            .in0(N__21975),
            .in1(N__16328),
            .in2(N__15834),
            .in3(N__19976),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_12_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_2_LC_9_8_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_2_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_2_LC_9_8_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_2_LC_9_8_4  (
            .in0(N__19247),
            .in1(N__15831),
            .in2(N__15819),
            .in3(N__19268),
            .lcout(\Lab_UT.scctrl.N_13_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNO_0_1_LC_9_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNO_0_1_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNO_0_1_LC_9_8_5 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \Lab_UT.scctrl.next_state_RNO_0_1_LC_9_8_5  (
            .in0(N__23180),
            .in1(N__18147),
            .in2(N__15816),
            .in3(N__16041),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_rst_0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_1_LC_9_8_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_1_LC_9_8_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.next_state_1_LC_9_8_6 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \Lab_UT.scctrl.next_state_1_LC_9_8_6  (
            .in0(N__16329),
            .in1(N__19977),
            .in2(N__16320),
            .in3(N__21976),
            .lcout(\Lab_UT.scctrl.next_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21119),
            .ce(N__20901),
            .sr(N__20846));
    defparam \Lab_UT.scctrl.state_2_fast_RNI7HMP_3_LC_9_9_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_fast_RNI7HMP_3_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_fast_RNI7HMP_3_LC_9_9_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \Lab_UT.scctrl.state_2_fast_RNI7HMP_3_LC_9_9_0  (
            .in0(N__16317),
            .in1(N__18898),
            .in2(_gnd_net_),
            .in3(N__16281),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_5_RNI7FV82_LC_9_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_5_RNI7FV82_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_5_RNI7FV82_LC_9_9_1 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_5_RNI7FV82_LC_9_9_1  (
            .in0(N__16163),
            .in1(N__16192),
            .in2(N__16257),
            .in3(N__16230),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_1_RNIGQ5R4_LC_9_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_1_RNIGQ5R4_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_1_RNIGQ5R4_LC_9_9_2 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_1_RNIGQ5R4_LC_9_9_2  (
            .in0(N__18247),
            .in1(N__16224),
            .in2(N__16254),
            .in3(N__23162),
            .lcout(\Lab_UT.scctrl.g0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_fast_RNIFRSV_2_LC_9_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_fast_RNIFRSV_2_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_fast_RNIFRSV_2_LC_9_9_3 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \Lab_UT.scctrl.state_1_fast_RNIFRSV_2_LC_9_9_3  (
            .in0(N__20375),
            .in1(N__21965),
            .in2(N__16164),
            .in3(N__16245),
            .lcout(\Lab_UT.scctrl.N_408_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_rep1_RNI9FBG_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNI9FBG_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_rep1_RNI9FBG_LC_9_9_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_rep1_RNI9FBG_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__19907),
            .in2(_gnd_net_),
            .in3(N__20512),
            .lcout(\Lab_UT.scctrl.g2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_19_LC_9_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_19_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_19_LC_9_9_5 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_19_LC_9_9_5  (
            .in0(N__20513),
            .in1(_gnd_net_),
            .in2(N__19934),
            .in3(N__18246),
            .lcout(\Lab_UT.scctrl.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_5_RNIH2CF_LC_9_9_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_5_RNIH2CF_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_5_RNIH2CF_LC_9_9_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_5_RNIH2CF_LC_9_9_6  (
            .in0(N__16191),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16162),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_412_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIJOFP1_LC_9_9_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIJOFP1_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNIJOFP1_LC_9_9_7 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNIJOFP1_LC_9_9_7  (
            .in0(N__18899),
            .in1(N__23573),
            .in2(N__16044),
            .in3(N__19596),
            .lcout(\Lab_UT.scctrl.next_state_rst_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_LC_9_10_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.nibbleIn1_LC_9_10_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_LC_9_10_0  (
            .in0(N__19749),
            .in1(N__16380),
            .in2(N__22593),
            .in3(N__16467),
            .lcout(\Lab_UT.scctrl.nibbleInZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21105),
            .ce(N__16497),
            .sr(N__16371));
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIQ5993_LC_9_10_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIQ5993_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIQ5993_LC_9_10_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_7_RNIQ5993_LC_9_10_1  (
            .in0(N__21972),
            .in1(N__22449),
            .in2(N__16485),
            .in3(N__22196),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_69_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNI6DT75_LC_9_10_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNI6DT75_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNI6DT75_LC_9_10_2 .LUT_INIT=16'b0000101000100010;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNI6DT75_LC_9_10_2  (
            .in0(N__21570),
            .in1(N__16466),
            .in2(N__16458),
            .in3(N__19748),
            .lcout(\Lab_UT.sccDnibble1En ),
            .ltout(\Lab_UT.sccDnibble1En_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_esr_RNO_2_LC_9_10_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_esr_RNO_2_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.u0.q_esr_RNO_2_LC_9_10_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.scdp.u0.q_esr_RNO_2_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16455),
            .in3(N__16452),
            .lcout(\Lab_UT.scdp.u0.sccDnibble1En_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIEAT93_LC_9_10_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIEAT93_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_7_RNIEAT93_LC_9_10_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_7_RNIEAT93_LC_9_10_4  (
            .in0(N__22198),
            .in1(N__16395),
            .in2(N__22463),
            .in3(N__21973),
            .lcout(\Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93 ),
            .ltout(\Lab_UT.scctrl.shifter_ret_7_RNIEATZ0Z93_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_0_LC_9_10_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_0_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_0_LC_9_10_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_0_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16374),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.scctrl.N_69_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_10_LC_9_10_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_10_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_10_LC_9_10_7 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_10_LC_9_10_7  (
            .in0(N__21971),
            .in1(N__22450),
            .in2(N__19031),
            .in3(N__22197),
            .lcout(\Lab_UT.scctrl.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIDAFVC_3_LC_9_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIDAFVC_3_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIDAFVC_3_LC_9_11_0 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIDAFVC_3_LC_9_11_0  (
            .in0(N__19620),
            .in1(N__23196),
            .in2(N__22977),
            .in3(N__16671),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_9_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIN96CP1_3_LC_9_11_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIN96CP1_3_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIN96CP1_3_LC_9_11_1 .LUT_INIT=16'b1100000000010000;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIN96CP1_3_LC_9_11_1  (
            .in0(N__16358),
            .in1(N__16716),
            .in2(N__16332),
            .in3(N__20017),
            .lcout(\Lab_UT.scctrl.next_state_RNIN96CP1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIV6006_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIV6006_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.shifter_ret_3_RNIV6006_LC_9_11_2 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \Lab_UT.scctrl.shifter_ret_3_RNIV6006_LC_9_11_2  (
            .in0(N__16755),
            .in1(N__16743),
            .in2(_gnd_net_),
            .in3(N__16730),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g1_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNICEBUC_3_LC_9_11_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNICEBUC_3_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNICEBUC_3_LC_9_11_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Lab_UT.scctrl.next_state_RNICEBUC_3_LC_9_11_3  (
            .in0(N__23454),
            .in1(N__19518),
            .in2(N__16719),
            .in3(N__16677),
            .lcout(\Lab_UT.scctrl.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNI91NK6_2_LC_9_11_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNI91NK6_2_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNI91NK6_2_LC_9_11_4 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNI91NK6_2_LC_9_11_4  (
            .in0(N__19103),
            .in1(N__16710),
            .in2(N__16704),
            .in3(N__23195),
            .lcout(\Lab_UT.scctrl.g0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIDJ6B1_2_LC_9_11_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIDJ6B1_2_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIDJ6B1_2_LC_9_11_5 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIDJ6B1_2_LC_9_11_5  (
            .in0(N__20313),
            .in1(N__19104),
            .in2(N__18429),
            .in3(N__22815),
            .lcout(\Lab_UT.scctrl.g0_9_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u1.q_3_LC_9_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_3_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u1.q_3_LC_9_12_0 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \Lab_UT.scdp.u1.q_3_LC_9_12_0  (
            .in0(N__21537),
            .in1(N__16661),
            .in2(N__17913),
            .in3(N__17893),
            .lcout(\Lab_UT.scdp.byteToDecrypt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21093),
            .ce(),
            .sr(N__20825));
    defparam \Lab_UT.scdp.a2b.val_i_0_0_LC_9_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_i_0_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_i_0_0_LC_9_12_1 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \Lab_UT.scdp.a2b.val_i_0_0_LC_9_12_1  (
            .in0(N__17055),
            .in1(N__16643),
            .in2(N__17206),
            .in3(N__17074),
            .lcout(\Lab_UT.scdp.val_i_0_0 ),
            .ltout(\Lab_UT.scdp.val_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.rxdataD.q_0_LC_9_12_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.rxdataD.q_0_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.rxdataD.q_0_LC_9_12_2 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \Lab_UT.scdp.rxdataD.q_0_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16647),
            .in3(N__17276),
            .lcout(\Lab_UT.scdp.binValD_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21093),
            .ce(),
            .sr(N__20825));
    defparam \Lab_UT.scdp.a2b.val_i_a2_0_LC_9_12_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.val_i_a2_0_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.val_i_a2_0_LC_9_12_3 .LUT_INIT=16'b0101000000010000;
    LogicCell40 \Lab_UT.scdp.a2b.val_i_a2_0_LC_9_12_3  (
            .in0(N__16644),
            .in1(N__17195),
            .in2(N__16581),
            .in3(N__17075),
            .lcout(\Lab_UT.scdp.N_378 ),
            .ltout(\Lab_UT.scdp.N_378_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_0_LC_9_12_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_0_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u0.q_0_LC_9_12_4 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \Lab_UT.scdp.u0.q_0_LC_9_12_4  (
            .in0(N__17291),
            .in1(N__17306),
            .in2(N__17313),
            .in3(N__16951),
            .lcout(\Lab_UT.scdp.byteToDecrypt_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21093),
            .ce(),
            .sr(N__20825));
    defparam \Lab_UT.scdp.u1.q_0_LC_9_12_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u1.q_0_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u1.q_0_LC_9_12_5 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \Lab_UT.scdp.u1.q_0_LC_9_12_5  (
            .in0(N__17292),
            .in1(N__17251),
            .in2(N__17280),
            .in3(N__21536),
            .lcout(\Lab_UT.scdp.u1.byteToDecryptZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21093),
            .ce(),
            .sr(N__20825));
    defparam \Lab_UT.scdp.a2b.shifter_ret_RNIJ2EC2_LC_9_12_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.a2b.shifter_ret_RNIJ2EC2_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scdp.a2b.shifter_ret_RNIJ2EC2_LC_9_12_6 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \Lab_UT.scdp.a2b.shifter_ret_RNIJ2EC2_LC_9_12_6  (
            .in0(N__17232),
            .in1(N__17191),
            .in2(N__17076),
            .in3(N__17054),
            .lcout(\Lab_UT.scdp.val_0_tz_3 ),
            .ltout(\Lab_UT.scdp.val_0_tz_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.u0.q_3_LC_9_12_7 .C_ON=1'b0;
    defparam \Lab_UT.scdp.u0.q_3_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.u0.q_3_LC_9_12_7 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \Lab_UT.scdp.u0.q_3_LC_9_12_7  (
            .in0(N__16952),
            .in1(N__16926),
            .in2(N__16932),
            .in3(N__17892),
            .lcout(\Lab_UT.scdp.byteToDecrypt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21093),
            .ce(),
            .sr(N__20825));
    defparam \Lab_UT.scdp.k2l.q_0_LC_9_13_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2l.q_0_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2l.q_0_LC_9_13_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.scdp.k2l.q_0_LC_9_13_0  (
            .in0(N__17600),
            .in1(N__18685),
            .in2(N__16907),
            .in3(N__17453),
            .lcout(\Lab_UT.scdp.key2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21088),
            .ce(),
            .sr(N__20828));
    defparam \Lab_UT.scdp.k2l.q_1_LC_9_13_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2l.q_1_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2l.q_1_LC_9_13_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.scdp.k2l.q_1_LC_9_13_1  (
            .in0(N__17454),
            .in1(N__18676),
            .in2(N__16886),
            .in3(N__17408),
            .lcout(\Lab_UT.scdp.key2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21088),
            .ce(),
            .sr(N__20828));
    defparam \Lab_UT.scdp.k3l.q_0_LC_9_13_2 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3l.q_0_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3l.q_0_LC_9_13_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.scdp.k3l.q_0_LC_9_13_2  (
            .in0(N__17601),
            .in1(N__18686),
            .in2(N__16868),
            .in3(N__17948),
            .lcout(\Lab_UT.scdp.key3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21088),
            .ce(),
            .sr(N__20828));
    defparam \Lab_UT.scdp.k3l.q_1_LC_9_13_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3l.q_1_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3l.q_1_LC_9_13_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.scdp.k3l.q_1_LC_9_13_3  (
            .in0(N__17949),
            .in1(N__18677),
            .in2(N__16844),
            .in3(N__17409),
            .lcout(\Lab_UT.scdp.key3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21088),
            .ce(),
            .sr(N__20828));
    defparam \Lab_UT.scdp.k3l.q_2_LC_9_13_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3l.q_2_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3l.q_2_LC_9_13_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k3l.q_2_LC_9_13_4  (
            .in0(N__18675),
            .in1(N__16826),
            .in2(N__16772),
            .in3(N__17950),
            .lcout(\Lab_UT.scdp.key3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21088),
            .ce(),
            .sr(N__20828));
    defparam \Lab_UT.scdp.k3l.q_3_LC_9_13_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k3l.q_3_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k3l.q_3_LC_9_13_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.scdp.k3l.q_3_LC_9_13_5  (
            .in0(N__17951),
            .in1(N__18678),
            .in2(N__17930),
            .in3(N__18517),
            .lcout(\Lab_UT.scdp.key3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21088),
            .ce(),
            .sr(N__20828));
    defparam \Lab_UT.scdp.rxdataD.q_3_LC_9_13_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.rxdataD.q_3_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.rxdataD.q_3_LC_9_13_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.scdp.rxdataD.q_3_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__17909),
            .in2(_gnd_net_),
            .in3(N__17886),
            .lcout(\Lab_UT.scdp.binValD_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21088),
            .ce(),
            .sr(N__20828));
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_9_13_7 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_9_13_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \buart.Z_rx.hh_RNIJ3K62_0_LC_9_13_7  (
            .in0(N__17792),
            .in1(N__17763),
            .in2(_gnd_net_),
            .in3(N__17734),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scdp.k0l.q_0_LC_9_14_0 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0l.q_0_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0l.q_0_LC_9_14_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k0l.q_0_LC_9_14_0  (
            .in0(N__18679),
            .in1(N__17615),
            .in2(N__17573),
            .in3(N__17544),
            .lcout(\Lab_UT.scdp.key0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21082),
            .ce(),
            .sr(N__20829));
    defparam \Lab_UT.scdp.k0l.q_1_LC_9_14_1 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k0l.q_1_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k0l.q_1_LC_9_14_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k0l.q_1_LC_9_14_1  (
            .in0(N__17545),
            .in1(N__17393),
            .in2(N__17525),
            .in3(N__18682),
            .lcout(\Lab_UT.scdp.key0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21082),
            .ce(),
            .sr(N__20829));
    defparam \Lab_UT.scdp.k1h.q_1_LC_9_14_3 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1h.q_1_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1h.q_1_LC_9_14_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k1h.q_1_LC_9_14_3  (
            .in0(N__18683),
            .in1(N__17394),
            .in2(N__17474),
            .in3(N__17504),
            .lcout(\Lab_UT.scdp.key1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21082),
            .ce(),
            .sr(N__20829));
    defparam \Lab_UT.scdp.k2l.q_3_LC_9_14_4 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2l.q_3_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2l.q_3_LC_9_14_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k2l.q_3_LC_9_14_4  (
            .in0(N__18681),
            .in1(N__18516),
            .in2(N__17426),
            .in3(N__17456),
            .lcout(\Lab_UT.scdp.key2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21082),
            .ce(),
            .sr(N__20829));
    defparam \Lab_UT.scdp.k1l.q_1_LC_9_14_5 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k1l.q_1_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k1l.q_1_LC_9_14_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k1l.q_1_LC_9_14_5  (
            .in0(N__18684),
            .in1(N__17395),
            .in2(N__17330),
            .in3(N__17357),
            .lcout(\Lab_UT.scdp.key1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21082),
            .ce(),
            .sr(N__20829));
    defparam \Lab_UT.scdp.k2h.q_3_LC_9_14_6 .C_ON=1'b0;
    defparam \Lab_UT.scdp.k2h.q_3_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scdp.k2h.q_3_LC_9_14_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.scdp.k2h.q_3_LC_9_14_6  (
            .in0(N__18680),
            .in1(N__18515),
            .in2(N__18458),
            .in3(N__18484),
            .lcout(\Lab_UT.scdp.key2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21082),
            .ce(),
            .sr(N__20829));
    defparam \Lab_UT.scctrl.next_state_RNO_1_1_LC_11_5_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNO_1_1_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNO_1_1_LC_11_5_0 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \Lab_UT.scctrl.next_state_RNO_1_1_LC_11_5_0  (
            .in0(N__18428),
            .in1(N__19930),
            .in2(_gnd_net_),
            .in3(N__18276),
            .lcout(\Lab_UT.scctrl.next_state_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_2_rep2_RNIB7181_LC_11_5_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_2_rep2_RNIB7181_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_2_rep2_RNIB7181_LC_11_5_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.scctrl.state_1_2_rep2_RNIB7181_LC_11_5_1  (
            .in0(N__22963),
            .in1(N__21961),
            .in2(_gnd_net_),
            .in3(N__18066),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIE6PO6_0_LC_11_5_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIE6PO6_0_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIE6PO6_0_LC_11_5_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIE6PO6_0_LC_11_5_2  (
            .in0(N__21416),
            .in1(N__22288),
            .in2(N__18132),
            .in3(N__21521),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIMNKBA_3_LC_11_5_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIMNKBA_3_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIMNKBA_3_LC_11_5_3 .LUT_INIT=16'b0000110000000100;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIMNKBA_3_LC_11_5_3  (
            .in0(N__22965),
            .in1(N__18129),
            .in2(N__18117),
            .in3(N__23188),
            .lcout(\Lab_UT.scctrl.next_state_rst_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_5_LC_11_5_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_5_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_0_RNO_5_LC_11_5_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_0_RNO_5_LC_11_5_4  (
            .in0(N__18067),
            .in1(_gnd_net_),
            .in2(N__22035),
            .in3(N__22964),
            .lcout(\Lab_UT.scctrl.N_319_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_10_LC_11_6_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_10_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_10_LC_11_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_10_LC_11_6_0  (
            .in0(N__19599),
            .in1(N__18072),
            .in2(_gnd_net_),
            .in3(N__21818),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_5_LC_11_6_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_5_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_5_LC_11_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_5_LC_11_6_1  (
            .in0(N__21403),
            .in1(N__23509),
            .in2(N__17955),
            .in3(N__21520),
            .lcout(\Lab_UT.scctrl.G_18_i_a9_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_4_LC_11_6_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_4_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_4_LC_11_6_2 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_4_LC_11_6_2  (
            .in0(N__19164),
            .in1(N__23182),
            .in2(N__23523),
            .in3(N__22957),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_18_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_0_LC_11_6_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_0_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_0_LC_11_6_3 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_0_LC_11_6_3  (
            .in0(N__18978),
            .in1(N__18972),
            .in2(N__18960),
            .in3(N__22291),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_18_i_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_LC_11_6_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_ret_9_LC_11_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_LC_11_6_4  (
            .in0(N__19188),
            .in1(N__19215),
            .in2(N__18957),
            .in3(N__20055),
            .lcout(\Lab_UT.scctrl.N_398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21139),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_10_LC_11_6_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_10_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_10_LC_11_6_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_10_LC_11_6_5  (
            .in0(N__21817),
            .in1(N__20434),
            .in2(_gnd_net_),
            .in3(N__19598),
            .lcout(\Lab_UT.scctrl.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNICEV81_LC_11_6_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNICEV81_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNICEV81_LC_11_6_6 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNICEV81_LC_11_6_6  (
            .in0(N__19935),
            .in1(N__21402),
            .in2(N__21949),
            .in3(N__20179),
            .lcout(\Lab_UT.scctrl.state_1_ret_1_RNICEVZ0Z81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNI8F771_LC_11_6_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNI8F771_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNI8F771_LC_11_6_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.scctrl.state_1_2_rep1_RNI8F771_LC_11_6_7  (
            .in0(N__21816),
            .in1(N__20433),
            .in2(_gnd_net_),
            .in3(N__19597),
            .lcout(\Lab_UT.scctrl.N_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_0_LC_11_7_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_0_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_4_RNO_0_LC_11_7_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_RNO_0_LC_11_7_0  (
            .in0(N__23506),
            .in1(N__18936),
            .in2(N__20288),
            .in3(N__18924),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_4_LC_11_7_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_4_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_ret_4_LC_11_7_1 .LUT_INIT=16'b1100110011001111;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_4_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__20181),
            .in2(N__18909),
            .in3(N__20053),
            .lcout(\Lab_UT.scctrl.N_260_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21131),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNO_1_0_LC_11_7_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNO_1_0_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNO_1_0_LC_11_7_2 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \Lab_UT.scctrl.state_1_RNO_1_0_LC_11_7_2  (
            .in0(N__18861),
            .in1(N__22830),
            .in2(N__18831),
            .in3(N__18812),
            .lcout(\Lab_UT.scctrl.g0_1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_1_LC_11_7_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_1_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_1_LC_11_7_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.scctrl.state_1_1_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__20180),
            .in2(_gnd_net_),
            .in3(N__20052),
            .lcout(\Lab_UT.scctrl.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21131),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_2_LC_11_7_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_2_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_2_LC_11_7_4 .LUT_INIT=16'b0010011110101111;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_2_LC_11_7_4  (
            .in0(N__23505),
            .in1(N__19272),
            .in2(N__20289),
            .in3(N__19251),
            .lcout(\Lab_UT.scctrl.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_6_LC_11_7_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_6_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_6_LC_11_7_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_6_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__23672),
            .in2(_gnd_net_),
            .in3(N__19519),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_1_LC_11_7_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_1_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_1_LC_11_7_6 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_1_LC_11_7_6  (
            .in0(N__19209),
            .in1(N__23504),
            .in2(N__19191),
            .in3(N__19390),
            .lcout(\Lab_UT.scctrl.N_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNO_9_LC_11_7_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_9_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNO_9_LC_11_7_7 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNO_9_LC_11_7_7  (
            .in0(N__22436),
            .in1(N__21872),
            .in2(N__19179),
            .in3(N__22287),
            .lcout(\Lab_UT.scctrl.N_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_11_LC_11_8_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_11_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.nibbleIn1_RNO_11_LC_11_8_0 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \Lab_UT.scctrl.nibbleIn1_RNO_11_LC_11_8_0  (
            .in0(N__22258),
            .in1(N__19133),
            .in2(N__19035),
            .in3(N__23178),
            .lcout(\Lab_UT.scctrl.N_21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_14_LC_11_8_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_14_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_14_LC_11_8_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_14_LC_11_8_1  (
            .in0(N__22432),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21854),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_10_i_o7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_7_LC_11_8_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_7_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_7_LC_11_8_2 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_7_LC_11_8_2  (
            .in0(N__22259),
            .in1(N__19727),
            .in2(N__18993),
            .in3(N__23508),
            .lcout(\Lab_UT.scctrl.N_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_0_LC_11_8_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_0_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_0_LC_11_8_3 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_0_LC_11_8_3  (
            .in0(N__21204),
            .in1(N__18990),
            .in2(N__22592),
            .in3(N__22260),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_24_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_LC_11_8_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.rst_ret_LC_11_8_4 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \Lab_UT.scctrl.rst_ret_LC_11_8_4  (
            .in0(N__22637),
            .in1(N__22470),
            .in2(N__19761),
            .in3(N__19758),
            .lcout(\Lab_UT.scctrl.rst_retZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21126),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_2_LC_11_8_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_2_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_0_RNIJFLD2_2_LC_11_8_5 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_RNIJFLD2_2_LC_11_8_5  (
            .in0(N__21858),
            .in1(N__19726),
            .in2(N__22458),
            .in3(N__22256),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_0_RNIUTK59_LC_11_8_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_0_RNIUTK59_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_0_RNIUTK59_LC_11_8_6 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \Lab_UT.scctrl.state_ret_0_RNIUTK59_LC_11_8_6  (
            .in0(N__22257),
            .in1(N__19542),
            .in2(N__19632),
            .in3(N__19629),
            .lcout(\Lab_UT.scctrl.g0_9_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNIV3EJ1_LC_11_8_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNIV3EJ1_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_2_rep1_RNIV3EJ1_LC_11_8_7 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \Lab_UT.scctrl.state_1_2_rep1_RNIV3EJ1_LC_11_8_7  (
            .in0(N__21404),
            .in1(N__19607),
            .in2(N__20457),
            .in3(N__21853),
            .lcout(\Lab_UT.scctrl.g0_9_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNIU5BF_4_LC_11_9_0 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNIU5BF_4_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNIU5BF_4_LC_11_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.reset_count_RNIU5BF_4_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__22582),
            .in2(_gnd_net_),
            .in3(N__23443),
            .lcout(N_21_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_18_LC_11_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_18_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_18_LC_11_9_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_18_LC_11_9_1  (
            .in0(N__19494),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20250),
            .lcout(),
            .ltout(\Lab_UT.scctrl.m90_i_o6_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_13_LC_11_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_13_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_13_LC_11_9_2 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_13_LC_11_9_2  (
            .in0(N__19433),
            .in1(N__22583),
            .in2(N__19410),
            .in3(N__23444),
            .lcout(\Lab_UT.scctrl.N_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_1_LC_11_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_1_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_1_LC_11_9_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_5_RNO_1_LC_11_9_3  (
            .in0(N__19407),
            .in1(N__19391),
            .in2(_gnd_net_),
            .in3(N__19341),
            .lcout(),
            .ltout(\Lab_UT.scctrl.g0_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_0_LC_11_9_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_0_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_5_RNO_0_LC_11_9_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_5_RNO_0_LC_11_9_4  (
            .in0(N__20252),
            .in1(N__23448),
            .in2(N__19287),
            .in3(N__19284),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_5_LC_11_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_5_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_ret_5_LC_11_9_5 .LUT_INIT=16'b1000100010001010;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_5_LC_11_9_5  (
            .in0(N__22584),
            .in1(N__20140),
            .in2(N__20331),
            .in3(N__20054),
            .lcout(\Lab_UT.scctrl.N_356_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21120),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_4_RNIDMQE_LC_11_9_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_4_RNIDMQE_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_4_RNIDMQE_LC_11_9_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_4_RNIDMQE_LC_11_9_6  (
            .in0(N__23604),
            .in1(N__20139),
            .in2(_gnd_net_),
            .in3(N__23442),
            .lcout(\Lab_UT.scctrl.g0_9_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_0_LC_11_9_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNO_0_LC_11_9_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNO_0_LC_11_9_7  (
            .in0(N__20301),
            .in1(N__20251),
            .in2(N__23502),
            .in3(N__20196),
            .lcout(\Lab_UT.scctrl.next_state_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_3_LC_11_10_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.scctrl.state_1_ret_3_LC_11_10_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_LC_11_10_0  (
            .in0(N__20182),
            .in1(N__20061),
            .in2(_gnd_net_),
            .in3(N__20045),
            .lcout(\Lab_UT.scctrl.N_260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21115),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_RNIFADO_0_LC_11_10_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_RNIFADO_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_RNIFADO_0_LC_11_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_RNIFADO_0_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__21413),
            .in2(_gnd_net_),
            .in3(N__21928),
            .lcout(),
            .ltout(\Lab_UT.scctrl.next_state_1_i_i_a2_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_ret_1_RNI4KSC6_LC_11_10_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNI4KSC6_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_1_RNI4KSC6_LC_11_10_2 .LUT_INIT=16'b1100110111111111;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_1_RNI4KSC6_LC_11_10_2  (
            .in0(N__19946),
            .in1(N__22194),
            .in2(N__19980),
            .in3(N__21518),
            .lcout(\Lab_UT.scctrl.next_state_rst_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNIP7S81_LC_11_10_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNIP7S81_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNIP7S81_LC_11_10_3 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNIP7S81_LC_11_10_3  (
            .in0(N__19956),
            .in1(N__21414),
            .in2(N__22030),
            .in3(N__19947),
            .lcout(N_74),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_RNIOCR32_LC_11_10_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_RNIOCR32_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_11_RNIOCR32_LC_11_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_RNIOCR32_LC_11_10_4  (
            .in0(N__22428),
            .in1(N__19815),
            .in2(N__19788),
            .in3(N__22193),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_72_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_11_RNI4RQC3_LC_11_10_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_11_RNI4RQC3_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_11_RNI4RQC3_LC_11_10_5 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \Lab_UT.scctrl.state_ret_11_RNI4RQC3_LC_11_10_5  (
            .in0(N__21187),
            .in1(N__19770),
            .in2(N__21627),
            .in3(N__21608),
            .lcout(\Lab_UT.state_ret_11_RNI4RQC3_0 ),
            .ltout(\Lab_UT.state_ret_11_RNI4RQC3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_9_RNIP7S81_0_LC_11_10_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_9_RNIP7S81_0_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_9_RNIP7S81_0_LC_11_10_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.scctrl.state_ret_9_RNIP7S81_0_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21597),
            .in3(N__21561),
            .lcout(\Lab_UT.sccDnibble2En ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_3_LC_11_10_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_3_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_3_LC_11_10_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_3_LC_11_10_7  (
            .in0(N__21519),
            .in1(N__21415),
            .in2(N__21219),
            .in3(N__23513),
            .lcout(\Lab_UT.scctrl.G_10_i_a7_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_2_LC_11_11_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_2_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.scctrl.next_state_2_LC_11_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.scctrl.next_state_2_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21188),
            .lcout(\Lab_UT.scctrl.next_state_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21107),
            .ce(N__20892),
            .sr(N__20858));
    defparam \Lab_UT.scctrl.state_1_ret_3_RNIJURV_LC_11_12_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNIJURV_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_ret_3_RNIJURV_LC_11_12_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.scctrl.state_1_ret_3_RNIJURV_LC_11_12_1  (
            .in0(N__20686),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20663),
            .lcout(N_55_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_17_LC_12_8_7 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_17_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_17_LC_12_8_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_17_LC_12_8_7  (
            .in0(N__20524),
            .in1(N__23503),
            .in2(N__20447),
            .in3(N__22821),
            .lcout(\Lab_UT.scctrl.N_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_11_LC_12_9_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_11_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_11_LC_12_9_0 .LUT_INIT=16'b1111111100110111;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_11_LC_12_9_0  (
            .in0(N__23440),
            .in1(N__23606),
            .in2(N__23695),
            .in3(N__20391),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_10_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_5_LC_12_9_1 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_5_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_5_LC_12_9_1 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_5_LC_12_9_1  (
            .in0(N__22962),
            .in1(N__23198),
            .in2(N__20385),
            .in3(N__23441),
            .lcout(\Lab_UT.scctrl.G_10_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_1_fast_RNIM0M4_2_LC_12_9_2 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_1_fast_RNIM0M4_2_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_1_fast_RNIM0M4_2_LC_12_9_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.scctrl.state_1_fast_RNIM0M4_2_LC_12_9_2  (
            .in0(N__20382),
            .in1(N__22788),
            .in2(N__23501),
            .in3(N__20358),
            .lcout(),
            .ltout(\Lab_UT.scctrl.N_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.next_state_RNIMPVR_2_LC_12_9_3 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.next_state_RNIMPVR_2_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.next_state_RNIMPVR_2_LC_12_9_3 .LUT_INIT=16'b1111001111110111;
    LogicCell40 \Lab_UT.scctrl.next_state_RNIMPVR_2_LC_12_9_3  (
            .in0(N__23668),
            .in1(N__23605),
            .in2(N__23532),
            .in3(N__23438),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_15_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_2_RNIKG4B3_3_LC_12_9_4 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_2_RNIKG4B3_3_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_2_RNIKG4B3_3_LC_12_9_4 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \Lab_UT.scctrl.state_2_RNIKG4B3_3_LC_12_9_4  (
            .in0(N__23439),
            .in1(N__23181),
            .in2(N__22980),
            .in3(N__22961),
            .lcout(\Lab_UT.scctrl.G_15_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_6_LC_12_9_5 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_6_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_6_LC_12_9_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_6_LC_12_9_5  (
            .in0(N__22789),
            .in1(N__22636),
            .in2(N__22617),
            .in3(N__21735),
            .lcout(),
            .ltout(\Lab_UT.scctrl.G_24_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_1_LC_12_9_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_1_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_1_LC_12_9_6 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_1_LC_12_9_6  (
            .in0(N__22608),
            .in1(N__22602),
            .in2(N__22596),
            .in3(N__22585),
            .lcout(\Lab_UT.scctrl.G_24_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.rst_ret_RNO_12_LC_12_10_6 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.rst_ret_RNO_12_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.rst_ret_RNO_12_LC_12_10_6 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \Lab_UT.scctrl.rst_ret_RNO_12_LC_12_10_6  (
            .in0(N__22459),
            .in1(N__22195),
            .in2(_gnd_net_),
            .in3(N__21948),
            .lcout(\Lab_UT.scctrl.N_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.scctrl.state_ret_13_RNICOE1_LC_12_12_0 .C_ON=1'b0;
    defparam \Lab_UT.scctrl.state_ret_13_RNICOE1_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.scctrl.state_ret_13_RNICOE1_LC_12_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.scctrl.state_ret_13_RNICOE1_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21722),
            .lcout(N_245_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // latticehx1k
